`ifndef ARCH_H
`define ARCH_H

// `define RV32I
`define RV64I
`define RVM
`define RVA
`define RVF
`define RVD
`define RVC
`define ZBA
`define ZBB
// `define DIFFTEST

`define EXT_FENCEI

`define FEAT_SC
`define FEAT_ITTAGE_REGION
`define FEAT_L2CACHE
`define FEAT_MEMPRED

// `define SYNTH_VIVADO

`include "predefine.svh"
`endif
