VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sky130_sram_1r1w0rw_11x512
   CLASS BLOCK ;
   SIZE 397.78 BY 392.53 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  75.6 0.0 75.98 0.38 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  81.44 0.0 81.82 0.38 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  87.28 0.0 87.66 0.38 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  93.12 0.0 93.5 0.38 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  98.96 0.0 99.34 0.38 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  104.8 0.0 105.18 0.38 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  110.64 0.0 111.02 0.38 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  116.48 0.0 116.86 0.38 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  122.32 0.0 122.7 0.38 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  128.16 0.0 128.54 0.38 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  134.0 0.0 134.38 0.38 ;
      END
   END din0[10]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  63.92 0.0 64.3 0.38 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  69.76 0.0 70.14 0.38 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 117.81 0.38 118.19 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 126.31 0.38 126.69 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 131.95 0.38 132.33 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 140.45 0.38 140.83 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 146.09 0.38 146.47 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 154.59 0.38 154.97 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 159.985 0.38 160.365 ;
      END
   END addr0[8]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  327.64 392.15 328.02 392.53 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  321.8 392.15 322.18 392.53 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  397.4 72.67 397.78 73.05 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  397.4 64.17 397.78 64.55 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  397.4 58.53 397.78 58.91 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  346.7 0.0 347.08 0.38 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  343.725 0.0 344.105 0.38 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  344.415 0.0 344.795 0.38 ;
      END
   END addr1[7]
   PIN addr1[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  345.16 0.0 345.54 0.38 ;
      END
   END addr1[8]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 24.0 0.38 24.38 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  397.4 372.46 397.78 372.84 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  30.26 0.0 30.64 0.38 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  367.14 392.15 367.52 392.53 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  130.485 392.15 130.865 392.53 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  142.965 392.15 143.345 392.53 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  155.445 392.15 155.825 392.53 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  167.925 392.15 168.305 392.53 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  180.405 392.15 180.785 392.53 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  192.885 392.15 193.265 392.53 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  205.365 392.15 205.745 392.53 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  217.845 392.15 218.225 392.53 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  230.325 392.15 230.705 392.53 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  242.805 392.15 243.185 392.53 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  255.285 392.15 255.665 392.53 ;
      END
   END dout1[10]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  0.0 0.0 1.74 392.53 ;
         LAYER met3 ;
         RECT  0.0 390.79 397.78 392.53 ;
         LAYER met3 ;
         RECT  0.0 0.0 397.78 1.74 ;
         LAYER met4 ;
         RECT  396.04 0.0 397.78 392.53 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  392.56 3.48 394.3 389.05 ;
         LAYER met3 ;
         RECT  3.48 387.31 394.3 389.05 ;
         LAYER met3 ;
         RECT  3.48 3.48 394.3 5.22 ;
         LAYER met4 ;
         RECT  3.48 3.48 5.22 389.05 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 397.16 391.91 ;
   LAYER  met2 ;
      RECT  0.62 0.62 397.16 391.91 ;
   LAYER  met3 ;
      RECT  0.98 117.21 397.16 118.79 ;
      RECT  0.62 118.79 0.98 125.71 ;
      RECT  0.62 127.29 0.98 131.35 ;
      RECT  0.62 132.93 0.98 139.85 ;
      RECT  0.62 141.43 0.98 145.49 ;
      RECT  0.62 147.07 0.98 153.99 ;
      RECT  0.62 155.57 0.98 159.385 ;
      RECT  0.98 72.07 396.8 73.65 ;
      RECT  0.98 73.65 396.8 117.21 ;
      RECT  396.8 73.65 397.16 117.21 ;
      RECT  396.8 65.15 397.16 72.07 ;
      RECT  396.8 59.51 397.16 63.57 ;
      RECT  0.62 24.98 0.98 117.21 ;
      RECT  0.98 118.79 396.8 371.86 ;
      RECT  0.98 371.86 396.8 373.44 ;
      RECT  396.8 118.79 397.16 371.86 ;
      RECT  0.62 160.965 0.98 390.19 ;
      RECT  396.8 373.44 397.16 390.19 ;
      RECT  396.8 2.34 397.16 57.93 ;
      RECT  0.62 2.34 0.98 23.4 ;
      RECT  0.98 373.44 2.88 386.71 ;
      RECT  0.98 386.71 2.88 389.65 ;
      RECT  0.98 389.65 2.88 390.19 ;
      RECT  2.88 373.44 394.9 386.71 ;
      RECT  2.88 389.65 394.9 390.19 ;
      RECT  394.9 373.44 396.8 386.71 ;
      RECT  394.9 386.71 396.8 389.65 ;
      RECT  394.9 389.65 396.8 390.19 ;
      RECT  0.98 2.34 2.88 2.88 ;
      RECT  0.98 2.88 2.88 5.82 ;
      RECT  0.98 5.82 2.88 72.07 ;
      RECT  2.88 2.34 394.9 2.88 ;
      RECT  2.88 5.82 394.9 72.07 ;
      RECT  394.9 2.34 396.8 2.88 ;
      RECT  394.9 2.88 396.8 5.82 ;
      RECT  394.9 5.82 396.8 72.07 ;
   LAYER  met4 ;
      RECT  75.0 0.98 76.58 391.91 ;
      RECT  76.58 0.62 80.84 0.98 ;
      RECT  82.42 0.62 86.68 0.98 ;
      RECT  88.26 0.62 92.52 0.98 ;
      RECT  94.1 0.62 98.36 0.98 ;
      RECT  99.94 0.62 104.2 0.98 ;
      RECT  105.78 0.62 110.04 0.98 ;
      RECT  111.62 0.62 115.88 0.98 ;
      RECT  117.46 0.62 121.72 0.98 ;
      RECT  123.3 0.62 127.56 0.98 ;
      RECT  129.14 0.62 133.4 0.98 ;
      RECT  64.9 0.62 69.16 0.98 ;
      RECT  70.74 0.62 75.0 0.98 ;
      RECT  76.58 0.98 327.04 391.55 ;
      RECT  327.04 0.98 328.62 391.55 ;
      RECT  322.78 391.55 327.04 391.91 ;
      RECT  134.98 0.62 343.125 0.98 ;
      RECT  31.24 0.62 63.32 0.98 ;
      RECT  328.62 391.55 366.54 391.91 ;
      RECT  76.58 391.55 129.885 391.91 ;
      RECT  131.465 391.55 142.365 391.91 ;
      RECT  143.945 391.55 154.845 391.91 ;
      RECT  156.425 391.55 167.325 391.91 ;
      RECT  168.905 391.55 179.805 391.91 ;
      RECT  181.385 391.55 192.285 391.91 ;
      RECT  193.865 391.55 204.765 391.91 ;
      RECT  206.345 391.55 217.245 391.91 ;
      RECT  218.825 391.55 229.725 391.91 ;
      RECT  231.305 391.55 242.205 391.91 ;
      RECT  243.785 391.55 254.685 391.91 ;
      RECT  256.265 391.55 321.2 391.91 ;
      RECT  2.34 0.62 29.66 0.98 ;
      RECT  347.68 0.62 395.44 0.98 ;
      RECT  368.12 391.55 395.44 391.91 ;
      RECT  328.62 0.98 391.96 2.88 ;
      RECT  328.62 2.88 391.96 389.65 ;
      RECT  328.62 389.65 391.96 391.55 ;
      RECT  391.96 0.98 394.9 2.88 ;
      RECT  391.96 389.65 394.9 391.55 ;
      RECT  394.9 0.98 395.44 2.88 ;
      RECT  394.9 2.88 395.44 389.65 ;
      RECT  394.9 389.65 395.44 391.55 ;
      RECT  2.34 0.98 2.88 2.88 ;
      RECT  2.34 2.88 2.88 389.65 ;
      RECT  2.34 389.65 2.88 391.91 ;
      RECT  2.88 0.98 5.82 2.88 ;
      RECT  2.88 389.65 5.82 391.91 ;
      RECT  5.82 0.98 75.0 2.88 ;
      RECT  5.82 2.88 75.0 389.65 ;
      RECT  5.82 389.65 75.0 391.91 ;
   END
END    sky130_sram_1r1w0rw_11x512
END    LIBRARY
