`ifndef DEFINES_SVH
`define DEFINES_SVH
`include "interfaces.svh"
`include "functions.svh"
`include "postdefine.svh"
`endif
