`include "../../defines/defines.svh"

// btb update: idx, updateEntry
// tage update: pred, pred error

module FSQ (
    input logic clk,
    input logic rst,
    BpuFsqIO.fsq bpu_fsq_io,
    FsqCacheIO.fsq fsq_cache_io,
    PreDecodeRedirect.redirect pd_redirect,
    FsqBackendIO.fsq fsq_back_io,
    CommitBus.in commitBus,
    input FrontendCtrl frontendCtrl
);
    // TODO: update branch predictor when squash. Because branch metas are stored in ram
    // so even Wrongly updated branch predictor, it can be recovered when update
    logic `N(`FSQ_WIDTH) search_head, commit_head, tail, write_index;
    logic `N(`FSQ_WIDTH) search_head_n1, tail_n1, n_commit_head;
    logic `N(`FSQ_WIDTH) write_tail;
    logic `N(`FSQ_WIDTH) squashIdx;
    logic full;
    logic queue_we;
    logic last_stage_we;
    logic cache_req;
    logic cache_req_ok;
    BTBUpdateInfo oldEntry, oldErrorEntry;
    logic `N(`FSQ_SIZE) directionTable;
    logic tdir, hdir, shdir;
    logic `N(`FSQ_WIDTH) searchIdx;
    FetchStream commitStream, searchStream, writeStream, redirectStream;
    logic `N(`PREDICTION_WIDTH) commitSize;
    logic initReady;
    logic commitValid;
    FetchStream `N(`ALU_SIZE) back_streams;
    BranchRedirectInfo rd_br;
    CSRRedirectInfo rd_csr;
    logic rd_br_en;
    logic `N(`FSQ_WIDTH) rd_br_idx;


    logic `N(`FSQ_WIDTH) exception_head, exception_head_n, exception_head_pre;
    logic `ARRAY(`COMMIT_WIDTH, `FSQ_WIDTH) commitFsqIdx;
    logic commit_exc_valid;
    logic `N(`COMMIT_WIDTH) commit_older;
    logic `N(`PREDICTION_WIDTH) pd_size;
    logic exc_wen;
    logic `N(`FSQ_WIDTH) exc_widx;
`ifdef RVC
    logic `N(`SLOT_NUM) exc_rvc_pre, exc_rvc, commit_slot_rvc;
    logic `N(`BLOCK_INST_SIZE) is_rvc, commit_is_rvc;
    logic commit_rd_rvc;
    logic `N(`BLOCK_INST_SIZE) commit_offset_dec, commit_offset_sel/*verilator split_var*/;
`endif
    logic `N(`VADDR_SIZE) exc_waddr;

    assign tail_n1 = tail + 1;
    assign search_head_n1 = search_head + 1;
    assign write_tail = bpu_fsq_io.redirect ? bpu_fsq_io.prediction.stream_idx : tail;
    assign queue_we = bpu_fsq_io.en & (~full | bpu_fsq_io.redirect);
    assign last_stage_we = bpu_fsq_io.lastStage & (~full | bpu_fsq_io.redirect);
    assign write_index = rd_br_en ? rd_br_idx :
                         pd_redirect.en ? pd_redirect.fsqIdx.idx :
                         bpu_fsq_io.redirect ? bpu_fsq_io.prediction.stream_idx : tail;
    assign searchIdx = fsq_back_io.redirect.en ? fsq_back_io.redirect.fsqInfo.idx : search_head;
    assign writeStream = rd_br_en ? redirectStream : 
                         pd_redirect.en ? pd_redirect.stream :
                            bpu_fsq_io.prediction.stream;
    // read ports: cache, wb, commit
    MPRAM #(
        .WIDTH($bits(FetchStream)),
        .DEPTH(`FSQ_SIZE),
        .READ_PORT(1 + `ALU_SIZE + 1),
        .WRITE_PORT(1),
        .RESET(1)
    ) fs_queue(
        .clk(clk),
        .rst(rst),
        .rst_sync(1'b0),
        .en({cache_req_ok | fsq_back_io.redirect.en, {(`ALU_SIZE+1){1'b1}}}),
        .we((queue_we | pd_redirect.en | rd_br_en)),
        .waddr(write_index),
        .raddr({searchIdx, fsq_back_io.fsqIdx, n_commit_head}),
        .wdata(writeStream),
        .rdata({searchStream, back_streams, commitStream}),
        .ready(initReady)
    );


    RedirectInfo u_redirectInfo, commit_redictInfo;
    assign squashIdx = rd_br.en | rd_csr.en ? fsq_back_io.redirect.fsqInfo.idx : pd_redirect.fsqIdx.idx;
    MPRAM #(
        .WIDTH($bits(RedirectInfo)),
        .DEPTH(`FSQ_SIZE),
        .READ_PORT(2),
        .WRITE_PORT(1),
        .RESET(1)
    ) redirect_ram (
        .clk(clk),
        .rst(rst),
        .rst_sync(1'b0),
        .en(2'b11),
        .we(bpu_fsq_io.lastStage),
        .waddr(bpu_fsq_io.lastStageIdx),
        .raddr({commit_head, squashIdx}),
        .wdata(bpu_fsq_io.lastStagePred.redirect_info),
        .rdata({commit_redictInfo, u_redirectInfo}),
        .ready()
    );

    wire pd_nobranch = pd_redirect.en & ~pd_redirect.direct;
    wire btb_we = queue_we | pd_nobranch;
    wire [`FSQ_WIDTH-1:0] btb_waddr = pd_nobranch ? pd_redirect.fsqIdx.idx : write_tail;
    MPRAM #(
        .WIDTH($bits(BTBUpdateInfo)),
        .DEPTH(`FSQ_SIZE),
        .READ_PORT(1),
        .WRITE_PORT(1),
        .RESET(1)
    ) btb_ram (
        .clk(clk),
        .rst(rst),
        .rst_sync(1'b0),
        .en(1'b1),
        .raddr(n_commit_head),
        .rdata(oldEntry),
        .we(btb_we),
        .waddr(btb_waddr),
        .wdata(pd_nobranch ? 0 : bpu_fsq_io.prediction.btbEntry),
        .ready()
    );

    PredictionMeta updateMeta;
    MPRAM #(
        .WIDTH($bits(PredictionMeta)),
        .DEPTH(`FSQ_SIZE),
        .READ_PORT(1),
        .WRITE_PORT(1),
        .RESET(1)
    ) meta_ram (
        .clk(clk),
        .rst(rst),
        .rst_sync(1'b0),
        .en(1'b1),
        .raddr(commit_head),
        .rdata(updateMeta),
        .we(bpu_fsq_io.lastStage),
        .waddr(bpu_fsq_io.lastStageIdx),
        .wdata(bpu_fsq_io.lastStageMeta),
        .ready()
    );

    // for predecode redirectdeocder_exccode
    MPRAM #(
        .WIDTH(`VADDR_SIZE),
        .DEPTH(`FSQ_SIZE),
        .READ_PORT(1),
        .WRITE_PORT(1)
    ) ras_addr_ram (
        .clk(clk),
        .rst(rst),
        .rst_sync(1'b0),
        .en(1'b1),
        .raddr(pd_redirect.fsqIdx_pre),
        .rdata(pd_redirect.ras_addr),
        .we(bpu_fsq_io.lastStage),
        .waddr(bpu_fsq_io.lastStageIdx),
        .wdata(bpu_fsq_io.ras_addr),
        .ready()
    );

    typedef struct packed {
        logic `N(2) condNum;
        logic `N(`SLOT_NUM) condHist;
        logic `N(`SLOT_NUM) condValid;
        logic `ARRAY(`SLOT_NUM, `PREDICTION_WIDTH) offsets;
    } PredictionInfo;

    PredictionInfo predictionInfos `N(`FSQ_SIZE);
    PredictionInfo pd_wr_info;
    logic `N(`SLOT_NUM) condSmallNum, pd_smallNum;
    logic `N(`SLOT_NUM) condSmallNumAll, pd_smallNumAll;
    logic redirectIsCond;
    PredictionInfo redirectPredInfo;
    PredictionInfo pd_predInfo;
    PredictionInfo u_predInfo;

    assign pd_wr_info.condNum = bpu_fsq_io.prediction.cond_num;
    assign pd_wr_info.condHist = bpu_fsq_io.prediction.predTaken;
    BTBUpdateInfo predEntry;
    assign predEntry = bpu_fsq_io.prediction.btbEntry;
generate
    for(genvar i=0; i<`SLOT_NUM-1; i++)begin
        assign pd_wr_info.offsets[i] = predEntry.slots[i].offset;
    end
    assign pd_wr_info.condValid = bpu_fsq_io.prediction.cond_valid;
    assign pd_wr_info.offsets[`SLOT_NUM-1] = predEntry.tailSlot.offset;
endgenerate

    always_ff @(posedge clk or negedge rst)begin
        if(rst == `RST)begin
            predictionInfos <= '{default: 0};
        end
        else begin
            if(btb_we)begin
                predictionInfos[btb_waddr] <= pd_nobranch ? 0 : pd_wr_info;
            end
        end
    end

// cache
    logic abandonStall;
    logic abandonStallCond;
    logic abandonStallPass;
    assign cache_req = ((search_head != tail) | (shdir ^ tdir)) & 
                       ~pd_redirect.en  & ~fsq_back_io.redirect.en;
    always_ff @(posedge clk)begin
        if(cache_req_ok | fsq_back_io.redirect.en | pd_redirect.en)begin
            fsq_cache_io.en <= cache_req;
            fsq_cache_io.fsqIdx.idx <= search_head;
            fsq_cache_io.fsqIdx.dir <= directionTable[search_head];
        end
        if(~((abandonStall | abandonStallCond) & (fsq_cache_io.stall | ~fsq_cache_io.ready)) | abandonStallPass)begin
            fsq_cache_io.abandon <= bpu_fsq_io.redirect;
            fsq_cache_io.abandonIdx.idx <= bpu_fsq_io.prediction.stream_idx;
            fsq_cache_io.abandonIdx.dir <= bpu_fsq_io.prediction.stream_dir;
            fsq_cache_io.abandonStream <= bpu_fsq_io.prediction.stream;
        end
    end

    assign abandonStallCond = fsq_cache_io.abandon & fsq_cache_io.abandonHit & (fsq_cache_io.stall | ~fsq_cache_io.ready);
    assign abandonStallPass = (abandonStall | abandonStallCond) & bpu_fsq_io.redirect & 
                            (fsq_cache_io.abandonIdx == {bpu_fsq_io.prediction.stream_idx, bpu_fsq_io.prediction.stream_dir});
    always_ff @(posedge clk or negedge rst)begin
        if(rst == `RST)begin
            abandonStall <= 1'b0;
        end
        else if(fsq_cache_io.flush)begin
            abandonStall <= 1'b0;
        end
        else begin
            if(abandonStallCond)begin
                abandonStall <= 1'b1;
            end
            else if(~fsq_cache_io.stall & fsq_cache_io.ready)begin
                abandonStall <= 1'b0;
            end
        end
    end
    assign fsq_cache_io.stream = searchStream;
    assign fsq_cache_io.flush = pd_redirect.en | fsq_back_io.redirect.en;
    assign fsq_cache_io.stall = frontendCtrl.ibuf_full;
    assign bpu_fsq_io.stream_idx = tail;
    assign bpu_fsq_io.stream_dir = tdir;
    assign bpu_fsq_io.stall = full;
    assign cache_req_ok = fsq_cache_io.ready;

    logic `N(`PREDICTION_WIDTH) shiftOffset, shiftIdx;
    always_ff @(posedge clk or negedge rst)begin
        if(rst == `RST)begin
            shiftOffset <= 0;
            shiftIdx <= 0;
        end
        else begin
            
            if(fsq_back_io.redirectBr.en | fsq_back_io.redirectCsr.en)begin
                shiftOffset <= 0;
                shiftIdx <= 0;
            end
            else if(fsq_back_io.redirect.en)begin
                // redirect mem, start from next instr
                shiftOffset <= fsq_back_io.redirect.fsqInfo.offset;
`ifdef RVC
                shiftIdx <= fsq_back_io.redirect.fsqInfo.size;
`endif
            end
            else if(cache_req_ok)begin
                shiftOffset <= 0;
                shiftIdx <= 0;
            end
        end
    end
    always_ff @(posedge clk)begin
        fsq_cache_io.shiftOffset <= shiftOffset;
`ifdef RVC
        fsq_cache_io.shiftIdx <= shiftIdx;
`endif
    end

    // logic `N(`SLOT_NUM) condFree;
    // PEncoder #(`SLOT_NUM) encoder_condFree({~oldEntry.slots[0].en, ~oldEntry.tailSlot.en}, condFree);

    CondPredInfo redirectCondInfo, pd_condInfo;
    assign pd_predInfo = predictionInfos[pd_redirect.fsqIdx.idx];
    assign redirectPredInfo = predictionInfos[fsq_back_io.redirect.fsqInfo.idx];

generate
    for(genvar i=0; i<`SLOT_NUM; i++)begin
        // 如果frontend redirect那么最后一个slot的类型一定不是cond
        assign pd_smallNum[i] = pd_predInfo.condValid[i] & (pd_predInfo.offsets[i] < pd_redirect.stream.size);
        assign condSmallNum[i] = redirectPredInfo.condValid[i] & (redirectPredInfo.offsets[i] < fsq_back_io.redirect.fsqInfo.offset);
    end
endgenerate
    assign redirectIsCond = fsq_back_io.redirectBr.en & fsq_back_io.redirectBr.br_type == CONDITION;
    `UNPARAM(SLOT_NUM, 2, "condSmallNum adder")
    assign condSmallNumAll = condSmallNum[0] + condSmallNum[1];
    wire [1:0] pd_smallMask;
    assign pd_smallMask[1] = pd_smallNum[1] & (&pd_smallNum);
    assign pd_smallMask[0] = pd_smallNum[0];
    assign pd_smallNumAll[1] = pd_smallMask[0] & pd_smallMask[1];
    assign pd_smallNumAll[0] = pd_smallMask[0] ^ pd_smallMask[1];
    
    assign pd_condInfo.condNum = {`SLOT_NUM{pd_redirect.stream.taken}} & pd_smallNumAll;
    assign pd_condInfo.taken = 0;
    always_comb begin
        if(redirectIsCond)begin
            if(condSmallNumAll < `SLOT_NUM)begin
                redirectCondInfo.condNum = condSmallNumAll + 1;
                redirectCondInfo.taken = fsq_back_io.redirectBr.taken;
            end
            else begin
                redirectCondInfo.condNum = `SLOT_NUM;
                redirectCondInfo.taken = 0;
            end
        end
        else begin
            redirectCondInfo.condNum = condSmallNumAll;
            redirectCondInfo.taken = 0;
        end
    end

// squash
    logic `N(`VADDR_SIZE) squash_target_pc;
    logic `N(`FSQ_WIDTH) pd_redirect_n1, bpu_fsq_redirect_n1, redirect_n1;
    logic rd_br_taken;
    logic `VADDR_BUS rd_br_target;
    logic `N(`PREDICTION_WIDTH) rd_br_offset;

    assign pd_redirect_n1 = pd_redirect.fsqIdx.idx + 1;
    assign bpu_fsq_redirect_n1 = bpu_fsq_io.prediction.stream_idx + 1;
    assign redirect_n1 = fsq_back_io.redirect.fsqInfo.idx + 1;

    CondPredInfo squash_pred_info;
    BranchType squash_br_type;
    logic squash_redirect_en, squash_pd_en;
    logic `VADDR_BUS pd_start_addr;
    logic `N(`PREDICTION_WIDTH) squash_offset;
    assign n_commit_head = commitValid ? commit_head + 1 : commit_head;
    assign full = commit_head == tail && (hdir ^ tdir);
    assign bpu_fsq_io.squashInfo.redirectInfo = u_redirectInfo;
    assign bpu_fsq_io.squashInfo.start_addr = squash_redirect_en ? searchStream.start_addr : pd_start_addr;
    assign bpu_fsq_io.squashInfo.offset = squash_offset;
    assign bpu_fsq_io.squashInfo.target_pc = squash_target_pc;
    assign bpu_fsq_io.squashInfo.predInfo = squash_pred_info;
    assign bpu_fsq_io.squashInfo.br_type = squash_br_type;
    assign bpu_fsq_io.squashInfo.squash_front = ~squash_redirect_en & squash_pd_en;
`ifdef DIFFTEST
    logic `N(`FSQ_WIDTH) squashIdx_n;
    `SIG_N(squashIdx, squashIdx_n)
    assign bpu_fsq_io.squashInfo.squashIdx = squashIdx_n;
`endif
    always_ff @(posedge clk)begin
        squash_redirect_en <= rd_br.en | rd_csr.en;
        squash_pd_en <= pd_redirect.en;
        pd_start_addr <= pd_redirect.stream.start_addr;
        bpu_fsq_io.squash <= pd_redirect.en | fsq_back_io.redirect.en & (rd_br.en | rd_csr.en);
        // bpu_fsq_io.squashInfo.redirectInfo <= u_redirectInfo;
        squash_target_pc <= rd_csr.en ? fsq_back_io.redirectCsr.exc_pc :
                            rd_br.en ? fsq_back_io.redirectBr.target : 
                                                        pd_redirect.stream.target;
        squash_pred_info <= rd_br.en | rd_csr.en ? redirectCondInfo : pd_condInfo;
        squash_br_type <= rd_br.en ? fsq_back_io.redirectBr.br_type : 
                          rd_csr.en ? DIRECT : pd_redirect.br_type;
        squash_offset <= rd_br.en | rd_csr.en ? fsq_back_io.redirect.fsqInfo.offset : pd_redirect.stream.size;
        rd_br_taken <= rd_br.taken;
        rd_br_target <= fsq_back_io.redirectBr.target;
        rd_br_offset <= fsq_back_io.redirect.fsqInfo.offset;
        rd_br_en <= fsq_back_io.redirect.en & rd_br.en;
        rd_br_idx <= fsq_back_io.redirect.fsqInfo.idx;
    end
    assign redirectStream.taken = rd_br_taken;
    assign redirectStream.start_addr = searchStream.start_addr;
    assign redirectStream.target = rd_br_target;
    assign redirectStream.size = rd_br_offset;
`ifdef RVC
    logic squash_rvc, rd_br_rvc;
    assign bpu_fsq_io.squashInfo.rvc = squash_rvc;
    assign redirectStream.rvc = rd_br_rvc;
    always_ff @(posedge clk)begin
        rd_br_rvc <= fsq_back_io.redirect.rvc;
        squash_rvc <= rd_br.en | rd_csr.en ? fsq_back_io.redirect.rvc : pd_redirect.stream.rvc;
    end
`endif

// idx maintain
    logic search_bigger, search_eq, search_abandon;
    LoopCompare #(`FSQ_WIDTH) cmp_redirect_search({bpu_fsq_io.prediction.stream_idx, bpu_fsq_io.prediction.stream_dir}, {search_head, shdir}, search_bigger);
    assign search_eq = {bpu_fsq_io.prediction.stream_idx, bpu_fsq_io.prediction.stream_dir} == {search_head, shdir};
    assign search_abandon = search_bigger;
    always_ff @(posedge clk or negedge rst)begin
        if(rst == `RST)begin
            search_head <= 0;
            commit_head <= 0;
            tail <= 0;
        end
        else begin
            if(fsq_back_io.redirectBr.en | fsq_back_io.redirectCsr.en)begin
                search_head <= redirect_n1;
            end
            else if(fsq_back_io.redirect.en)begin
                search_head <= fsq_back_io.redirect.fsqInfo.idx;
            end
            else if(pd_redirect.en)begin
                if(pd_redirect.direct)begin
                    search_head <= pd_redirect_n1;
                end
                else begin
                    search_head <= pd_redirect.fsqIdx.idx;
                end
            end
            else if(bpu_fsq_io.redirect & search_abandon)begin
                search_head <= bpu_fsq_redirect_n1;
            end
            else if(cache_req_ok & cache_req) begin
                search_head <= search_head_n1;
            end

            if(fsq_back_io.redirect.en & (rd_br.en | rd_csr.en))begin
                tail <= redirect_n1;
            end
            else if(pd_redirect.en)begin
                tail <= pd_redirect_n1;
            end
            else if(bpu_fsq_io.redirect)begin
                tail <= bpu_fsq_redirect_n1;
            end
            else if(bpu_fsq_io.en & ~full)begin
                tail <= tail_n1;
            end

            commit_head <= n_commit_head;
        end
    end

    logic `N(`FSQ_WIDTH) redirect_dir_idx, redirect_dir_idx_n1;
    assign redirect_dir_idx = fsq_back_io.redirect.fsqInfo.idx;

    always_ff @(posedge clk or negedge rst)begin
        if(rst == `RST)begin
            tdir <= 0;
            hdir <= 0;
            shdir <= 0;
            directionTable <= '{default: 0};
        end
        else begin
            if(fsq_back_io.redirect.en & (rd_br.en | rd_csr.en))begin
                tdir <= redirect_dir_idx[`FSQ_WIDTH-1] & ~redirect_n1[`FSQ_WIDTH-1] ? ~directionTable[redirect_dir_idx] : directionTable[redirect_dir_idx];
            end
            else if(pd_redirect.en)begin
                tdir <= pd_redirect.fsqIdx.idx[`FSQ_WIDTH-1] & ~pd_redirect_n1[`FSQ_WIDTH-1] ? ~pd_redirect.fsqIdx.dir : pd_redirect.fsqIdx.dir;
            end
            else if(bpu_fsq_io.redirect)begin
                tdir <= bpu_fsq_io.prediction.stream_idx[`FSQ_WIDTH-1] & ~bpu_fsq_redirect_n1[`FSQ_WIDTH-1] ? ~bpu_fsq_io.prediction.stream_dir : bpu_fsq_io.prediction.stream_dir;
            end
            else if(bpu_fsq_io.en & ~full)begin
                tdir <= tail[`FSQ_WIDTH-1] & ~tail_n1[`FSQ_WIDTH-1] ? ~tdir : tdir;
            end

            if(fsq_back_io.redirectBr.en | fsq_back_io.redirectCsr.en)begin
                shdir <= redirect_dir_idx[`FSQ_WIDTH-1] & ~redirect_n1[`FSQ_WIDTH-1] ? ~directionTable[redirect_dir_idx] : directionTable[redirect_dir_idx];
            end
            else if(fsq_back_io.redirect.en)begin
                shdir <= directionTable[redirect_dir_idx];
            end
            else if(pd_redirect.en)begin
                if(pd_redirect.direct)begin
                    shdir <= pd_redirect.fsqIdx.idx[`FSQ_WIDTH-1] & ~pd_redirect_n1[`FSQ_WIDTH-1] ? ~pd_redirect.fsqIdx.dir : pd_redirect.fsqIdx.dir;
                end
                else begin
                    shdir <= pd_redirect.fsqIdx.dir;
                end
            end
            else if(bpu_fsq_io.redirect & search_abandon)begin
                shdir <= bpu_fsq_io.prediction.stream_idx[`FSQ_WIDTH-1] & ~bpu_fsq_redirect_n1[`FSQ_WIDTH-1] ? ~bpu_fsq_io.prediction.stream_dir : bpu_fsq_io.prediction.stream_dir;
            end
            else if(cache_req_ok & cache_req)begin
                shdir <= search_head[`FSQ_WIDTH-1] & ~search_head_n1[`FSQ_WIDTH-1] ? ~shdir : shdir;
            end

            if(commitValid)begin
                hdir <= commit_head[`FSQ_WIDTH-1] & ~n_commit_head[`FSQ_WIDTH-1] ? ~hdir : hdir;
            end

            if(bpu_fsq_io.en & ~full)begin
                directionTable[tail] <= tdir;
            end
        end
    end

// wb & commit
    typedef struct packed {
`ifdef DIFFTEST
        logic front;
`endif
        logic exception;
        logic taken;
`ifdef RVC
        logic rvc;
        logic `N(`PREDICTION_WIDTH) size;
`endif
        BranchType br_type;
        logic `N(`VADDR_SIZE) target;
        logic `N(`PREDICTION_WIDTH) offset;
    } WBInfo;

    WBInfo wbInfos `N(`FSQ_SIZE);
    WBInfo commitWBInfo;
    logic `N(`FSQ_SIZE) pred_error_en, entry_error;
    logic pred_error;

    assign rd_br = fsq_back_io.redirectBr;
    assign rd_csr = fsq_back_io.redirectCsr;
    always_ff @(posedge clk or negedge rst)begin
        if(rst == `RST)begin
            wbInfos <= '{default: 0};
            pred_error_en <= 0;
            entry_error <= 0;
        end
        else begin
            if(pd_redirect.en)begin
                wbInfos[pd_redirect.fsqIdx.idx] <= {
`ifdef DIFFTEST
                1'b1,
`endif    
                1'b0, pd_redirect.direct,
`ifdef RVC
                pd_redirect.stream.rvc, pd_redirect.size,
`endif
                pd_redirect.br_type, 
                pd_redirect.stream.target, pd_redirect.stream.size};
            end
            if(rd_br.en | rd_csr.en)begin
                wbInfos[fsq_back_io.redirect.fsqInfo.idx] <= {
`ifdef DIFFTEST
                1'b0,
`endif
                rd_csr.en, rd_br.taken, 
`ifdef RVC
                fsq_back_io.redirect.rvc, fsq_back_io.redirect.fsqInfo.size,
`endif
                rd_br.br_type, rd_br.target, fsq_back_io.redirect.fsqInfo.offset};
            end
            if(queue_we)begin
                pred_error_en[write_index] <= 1'b0;
            end
            if(fsq_back_io.redirect.en & (rd_br.en | rd_csr.en))begin
                pred_error_en[fsq_back_io.redirect.fsqInfo.idx] <= 1'b1;
            end
            if(pd_redirect.en & pd_redirect.direct)begin
                pred_error_en[pd_redirect.fsqIdx.idx] <= 1'b1;
            end
            if(queue_we)begin
                entry_error[write_index] <= 1'b0;
            end
            if(pd_redirect.en & pd_redirect.entry_error)begin
                entry_error[pd_redirect.fsqIdx.idx] <= 1'b1;
            end
        end
    end

    localparam FSQ_INST_WIDTH=$clog2(`FSQ_SIZE*`BLOCK_INST_SIZE);
    logic `N(FSQ_INST_WIDTH+1) commitNum;
    BTBUpdateInfo commitUpdateEntry;
    FsqIdxInfo commitFsqInfo;
    logic `N(`PREDICTION_WIDTH) commitFsqSize;
`ifdef RVC
    assign commitFsqSize = commitWBInfo.size;
`else
    assign commitFsqSize = commitWBInfo.offset;
`endif
    // because streamVec is not init
    assign commitValid = initReady & (
                        (|commitNum[FSQ_INST_WIDTH: `PREDICTION_WIDTH]) || 
                        (commitNum[`PREDICTION_WIDTH-1: 0] > commitSize) ||
                        (pred_error_en[commit_head] & (commitNum[`PREDICTION_WIDTH-1: 0] > commitFsqSize)));
    assign pred_error = initReady & pred_error_en[commit_head] & 
                        ((|commitNum[FSQ_INST_WIDTH: `PREDICTION_WIDTH]) | (commitNum[`PREDICTION_WIDTH-1: 0] > commitFsqSize));

    logic `N(`PREDICTION_WIDTH) streamCommitSize;
    logic `N(`PREDICTION_WIDTH+1) streamCommitNum;

    assign streamCommitSize = pred_error_en[commit_head] ? commitFsqSize : commitSize;
    assign streamCommitNum = streamCommitSize + 1;

    always_ff @(posedge clk or negedge rst)begin
        if(rst == `RST)begin
            commitNum <= 0;
        end
        else begin
            commitNum <= commitNum + commitBus.num - ({`PREDICTION_WIDTH+1{commitValid}} & streamCommitNum);
        end
    end

    logic `N(`SLOT_NUM) realTaken, allocSlot;
    assign commitWBInfo = wbInfos[commit_head];
    assign u_predInfo = predictionInfos[commitFsqInfo.idx];
    assign commitFsqInfo.idx = commit_head;
`ifdef RVC
    assign commitFsqInfo.size = commitWBInfo.size;
`endif
    assign commitFsqInfo.offset = commitWBInfo.offset;
    assign oldErrorEntry = entry_error[commit_head] ? 0 : oldEntry;
    BTBEntryGen commit_btb_entry_gen (
        .oldEntry(oldErrorEntry),
        .pc(commitStream.start_addr),
        .fsqInfo(commitFsqInfo),
        .normalOffset(commitStream.size),
        .br_type(commitWBInfo.br_type),
        .pred_error(pred_error),
        .exception(commitWBInfo.exception),
        .target(commitWBInfo.target),
        .taken(commitWBInfo.taken),
`ifdef RVC
        .rvc(commitWBInfo.rvc),
        .slot_rvc(commit_slot_rvc),
        .rd_rvc(commit_rd_rvc),
`endif
        .predTaken(u_predInfo.condHist),
        .updateEntry(commitUpdateEntry),
        .realTaken(realTaken),
        .allocSlot(allocSlot)
    );

    logic update_taken, update_tail_taken;
    logic `N(`VADDR_SIZE) update_start_addr;
    logic `N(`VADDR_SIZE) update_target_pc, update_target_pc_pre;
    BTBUpdateInfo update_btb_entry, update_btb_entry_pre;
    PredErrorInfo update_error_info_pre, update_error_info;
    logic update_indirect, btb_update;
    logic `N(`SLOT_NUM) update_real_taken;
    logic `N(`SLOT_NUM) update_alloc_slot;
    assign bpu_fsq_io.updateInfo.meta = updateMeta;
    assign bpu_fsq_io.updateInfo.taken = update_taken;
    assign bpu_fsq_io.updateInfo.start_addr = update_start_addr;
    assign bpu_fsq_io.updateInfo.target_pc = update_target_pc;
    assign bpu_fsq_io.updateInfo.btbEntry = update_btb_entry;
    assign bpu_fsq_io.updateInfo.realTaken = update_real_taken;
    assign bpu_fsq_io.updateInfo.allocSlot = update_alloc_slot;
    assign bpu_fsq_io.updateInfo.tailTaken = update_tail_taken;
    assign bpu_fsq_io.updateInfo.redirectInfo = commit_redictInfo;
    assign bpu_fsq_io.updateInfo.btb_update = btb_update;
    assign bpu_fsq_io.updateInfo.error_info = update_error_info;
`ifdef DIFFTEST
    logic `N(`FSQ_WIDTH) dbg_commit_head;
    `SIG_N(commit_head, dbg_commit_head)
    assign bpu_fsq_io.updateInfo.fsqIdx = dbg_commit_head;
`endif
    assign update_target_pc_pre = pred_error ? commitWBInfo.target : commitStream.target;
`ifdef FEAT_ITTAGE_REGION
    assign bpu_fsq_io.ittage_tag = update_target_pc_pre[`ITTAGE_OFFSET + 1 +: `ITTAGE_REGION_TAG];
`endif
    assign update_error_info_pre.pred_error = pred_error;
    assign update_error_info_pre.fsqInfo = commitFsqInfo;
    assign update_error_info_pre.br_type = commitWBInfo.br_type;
`ifdef RVC
    assign update_error_info_pre.rvc = commitWBInfo.rvc;
`endif
    always_ff @(posedge clk)begin
        bpu_fsq_io.update <= commitValid;
        update_taken <= commitWBInfo.taken;
        update_start_addr <= commitStream.start_addr;
        update_target_pc <= update_target_pc_pre;
        update_btb_entry_pre <= pred_error ? commitUpdateEntry : oldErrorEntry;
        btb_update <= entry_error[commit_head] | pred_error & commitUpdateEntry.en;
        update_real_taken <= realTaken;
        update_alloc_slot <= allocSlot;
        update_tail_taken <= pred_error ? (commitWBInfo.br_type != CONDITION) & ~commitWBInfo.exception :
                            ~(|u_predInfo.condHist) & commitStream.taken;
        update_indirect <= pred_error ? commitWBInfo.br_type == INDIRECT || commitWBInfo.br_type == INDIRECT_CALL : 
                            ~(|u_predInfo.condHist) & commitStream.taken & ((oldEntry.tailSlot.br_type == INDIRECT) | (oldEntry.tailSlot.br_type == INDIRECT_CALL));
        update_error_info <= update_error_info_pre;
    end
    always_comb begin
        update_btb_entry = update_btb_entry_pre;
`ifdef FEAT_ITTAGE_REGION
        if(update_indirect)begin
            update_btb_entry.tailSlot.target[`ITTAGE_REGION_WIDTH-1: 0] = bpu_fsq_io.ittage_idx; 
        end
`endif
    end


generate
    for(genvar i=0; i<`COMMIT_WIDTH; i++)begin
        assign commit_older[i] = commitBus.en[i] & (commitBus.fsqInfo[i].idx != exception_head);
        assign commitFsqIdx[i] = commitBus.fsqInfo[i].idx;
    end
`ifdef RVC
    // 判断当前指令的前一条指令是否为rvc
    // 只需要前面两个槽，如果是rvi指令，那么前面两个槽都被占用
    // 则前面两个槽都不是rvc
    for(genvar i=0; i<`SLOT_NUM; i++)begin
        logic `N(`BLOCK_INST_SIZE) offset_dec;
        logic `N(`BLOCK_INST_SIZE) offset_sel/*verilator split_var*/;
        Decoder #(`BLOCK_INST_SIZE) decoder_br_offset (pd_predInfo.offsets[i], offset_dec);
        for(genvar j=0; j<`BLOCK_INST_SIZE-2; j++)begin
            assign offset_sel[j] = offset_dec[j+1] | offset_dec[j+2];
        end
        assign offset_sel[`BLOCK_INST_SIZE-2] = offset_dec[`BLOCK_INST_SIZE-1];
        assign offset_sel[`BLOCK_INST_SIZE-1] = 1'b0;
        wire `N(`BLOCK_INST_SIZE) rvc_mask = pd_redirect.is_rvc & offset_sel;
        assign exc_rvc_pre[i] = |rvc_mask;
    end
    Decoder #(`BLOCK_INST_SIZE) decoder_commit_offset (commitFsqInfo.offset, commit_offset_dec);
    for(genvar i=0; i<`BLOCK_INST_SIZE-2; i++)begin
        assign commit_offset_sel[i] = commit_offset_dec[i+1] | commit_offset_dec[i+2];
    end
    assign commit_offset_sel[`BLOCK_INST_SIZE-2] = commit_offset_dec[`BLOCK_INST_SIZE-1];
    assign commit_offset_sel[`BLOCK_INST_SIZE-1] = 1'b0;
    assign commit_rd_rvc = |(commit_offset_sel & commit_is_rvc);
`endif
endgenerate
    OldestSelect #(`COMMIT_WIDTH, 1, `FSQ_WIDTH) select_exception_head (
        commit_older, commitFsqIdx, commit_exc_valid, exception_head_n
    );
    always_ff @(posedge clk)begin
        exc_wen <= pd_redirect.exc_en;
        exc_widx <= pd_redirect.fsqIdx.idx;
        exc_waddr <= pd_redirect.stream.start_addr;
`ifdef RVC
        exc_rvc <= exc_rvc_pre;
        is_rvc <= pd_redirect.is_rvc;
`endif
        pd_size <= pd_redirect.size;
        exception_head_pre <= exception_head;
    end
    always_ff @(posedge clk, negedge rst)begin
        if(rst == `RST)begin
            exception_head <= 0;
        end
        else begin
            if(commit_exc_valid)begin
                exception_head <= exception_head_n;
            end
        end
    end

    logic `ARRAY(`COMMIT_WIDTH, `FSQ_WIDTH) exception_idxs;
    logic `ARRAY(`COMMIT_WIDTH, `PREDICTION_WIDTH+`VADDR_SIZE) exception_addrs;
generate
    for(genvar i=0; i<`COMMIT_WIDTH; i++)begin
        assign exception_idxs[i] = exception_head + i;
    end
endgenerate
    MPRAM #(
        .WIDTH(`VADDR_SIZE+`PREDICTION_WIDTH),
        .DEPTH(`FSQ_SIZE),
        .READ_PORT(`COMMIT_WIDTH),
        .WRITE_PORT(1)
    ) exception_ram (
        .clk(clk),
        .rst(rst),
        .rst_sync(1'b0),
        .en({`COMMIT_WIDTH{1'b1}}),
        .raddr(exception_idxs),
        .rdata(exception_addrs),
        .we(exc_wen),
        .waddr(exc_widx),
        .wdata({pd_size, exc_waddr}),
        .ready()
    );
    MPRAM #(
        .WIDTH(`PREDICTION_WIDTH
        `ifdef RVC
        +`SLOT_NUM + `BLOCK_INST_SIZE
        `endif),
        .DEPTH(`FSQ_SIZE),
        .READ_PORT(1),
        .WRITE_PORT(1)
    ) stream_size_ram (
        .clk(clk),
        .rst(rst),
        .rst_sync(1'b0),
        .en(1'b1),
        .raddr(n_commit_head),
        .rdata({commitSize
        `ifdef RVC
        ,{commit_slot_rvc, commit_is_rvc}
        `endif
        }),
        .we(exc_wen),
        .waddr(exc_widx),
        .wdata({pd_size
        `ifdef RVC
        ,{exc_rvc, is_rvc}
        `endif
        }),
        .ready()
    );
    logic `N($clog2(`COMMIT_WIDTH)) exc_stream_idx;
    assign exc_stream_idx = commitBus.fsqInfo[0].idx - exception_head_pre;
    assign fsq_back_io.commitStreamSize = exception_addrs[exc_stream_idx][`VADDR_SIZE +: `PREDICTION_WIDTH];

`ifdef RVC
    logic `N(`FSQ_SIZE) commit_head_mask, redirect_mask;
    logic `ARRAY(`ALU_SIZE, `PREDICTION_WIDTH) stream_lasts;
    logic `N(`PREDICTION_WIDTH) last_offset;
    always_ff @(posedge clk)begin
        last_offset <= pd_redirect.last_offset;
    end
    MaskGen #(`FSQ_SIZE) mask_gen_commit_head (commit_head, commit_head_mask);
    MaskGen #(`FSQ_SIZE) mask_gen_redirect (fsq_back_io.redirect.fsqInfo.idx, redirect_mask);

    MPRAM #(
        .WIDTH(`PREDICTION_WIDTH),
        .DEPTH(`FSQ_SIZE),
        .READ_PORT(`ALU_SIZE),
        .WRITE_PORT(1)
    ) stream_last_ram (
        .clk(clk),
        .rst(rst),
        .rst_sync(1'b0),
        .en({`ALU_SIZE{1'b1}}),
        .raddr(fsq_back_io.fsqIdx),
        .rdata(stream_lasts),
        .we(exc_wen),
        .waddr(exc_widx),
        .wdata(last_offset),
        .ready()
    );
generate
    for(genvar i=0; i<`ALU_SIZE; i++)begin
        always_comb begin
            fsq_back_io.streams[i] = back_streams[i];
            fsq_back_io.streams[i].size = stream_lasts[i];
        end
    end
endgenerate
`else
    assign fsq_back_io.streams = back_streams;
`endif

    logic `N($clog2(`COMMIT_WIDTH)) exc_ridx;
    assign exc_ridx = fsq_back_io.redirect.fsqInfo.idx - exception_head_pre;
    assign fsq_back_io.exc_pc = exception_addrs[exc_ridx][`VADDR_SIZE-1: 0] + {fsq_back_io.redirect.fsqInfo.offset, {`INST_OFFSET{1'b0}}};

`ifdef DIFFTEST
    logic `N(`VADDR_SIZE) diff_pcs `N(`FSQ_SIZE);
generate
    for(genvar i=0; i<`COMMIT_WIDTH; i++)begin
        assign fsq_back_io.diff_pc[i] = diff_pcs[fsq_back_io.diff_fsqInfo[i].idx] + {fsq_back_io.diff_fsqInfo[i].offset, {`INST_OFFSET{1'b0}}};
    end
endgenerate
    always_ff @(posedge clk or negedge rst)begin
        if(rst == `RST)begin
            diff_pcs <= '{default: 0};
        end
        else begin
            if(queue_we)begin
                diff_pcs[write_tail] <= bpu_fsq_io.prediction.stream.start_addr;
            end
            
        end
    end
    FetchStream logStream;
    logic logError;
    logic redirect_n;
    logic `N(`FSQ_WIDTH) redirect_idx;
    always_ff @(posedge clk)begin
        logStream <= commitStream;
        logError <= pred_error;
        redirect_n <= fsq_back_io.redirect.en;
        redirect_idx <= fsq_back_io.redirect.fsqInfo.idx;
    end
    `Log(DLog::Debug, T_FSQ, bpu_fsq_io.update, $sformatf("update BP%4d. [%8h %4d]->%8h %8h %b", commit_head, logStream.start_addr, logStream.size, logStream.target, update_target_pc, logError))
    `Log(DLog::Debug, T_FSQ, bpu_fsq_io.squash, $sformatf("squash BP [%d %d].", redirect_idx, redirect_n))

    `PERF(pred_error_cond, commitValid & pred_error & ~commitWBInfo.exception & commitWBInfo.br_type == CONDITION)
    `PERF(pred_error_ind, commitValid & pred_error & ~commitWBInfo.exception & 
    ((commitWBInfo.br_type == INDIRECT) | (commitWBInfo.br_type == INDIRECT_CALL)))
    `PERF(pred_error_call, commitValid & pred_error & ~commitWBInfo.exception & ~commitWBInfo.front & 
    ((commitWBInfo.br_type == POP) | (commitWBInfo.br_type == POP_PUSH) | (commitWBInfo.br_type == PUSH)))
    `PERF(pred_error, commitValid & pred_error & ~commitWBInfo.exception & ~commitWBInfo.front)
    `PERF(front_redirect_direct, pd_redirect.en & pd_redirect.direct)
    `PERF(front_redirect_nobranch, pd_redirect.en & ~pd_redirect.direct)

//     logic `N(6) dbg_commit_idx, dbg_commit_head;
//     logic `ARRAY(64, `FSQ_WIDTH) dbg_fsq_idxs;
//     logic `ARRAY(`COMMIT_WIDTH, 6) dbg_commit_idxs;
//     logic `ARRAY(8, 6) dbg_commit_head_idxs;

// generate
//     for(genvar i=0; i<`COMMIT_WIDTH; i++)begin
//         assign dbg_commit_idxs[i] = dbg_commit_idx + i;
//     end
//     for(genvar i=0; i<8; i++)begin
//         assign dbg_commit_head_idxs[i] = dbg_commit_head + i;
//     end
// endgenerate

//     always_ff @(posedge clk, negedge rst)begin
//         if(rst == `RST)begin
//             dbg_commit_idx <= 0;
//             dbg_fsq_idxs <= 0;
//             dbg_commit_head <= 0;
//         end
//         else begin
//             if(commitValid)begin
//                 dbg_commit_head <= dbg_commit_head + streamCommitNum;
//             end
//             dbg_commit_idx <= dbg_commit_idx + commitBus.num;
//             for(int i=0; i<`COMMIT_WIDTH; i++)begin
//                 if(i < commitBus.num)begin
//                     dbg_fsq_idxs[dbg_commit_idxs[i]] <= commitBus.fsqInfo[i].idx;
//                 end
//             end
//         end
//     end

//     always_ff @(posedge clk)begin
//         if(commitValid)begin
//             for(int i=0; i<8; i++)begin
//                 if((i < streamCommitNum) && commit_head != dbg_fsq_idxs[dbg_commit_head_idxs[i]])begin
//                     $display("[%16d] fsq commit[%d] error", DLog::cycleCnt, commit_head);
//                 end
//             end
//         end
//     end
`endif

endmodule

module BTBEntryGen(
    input BTBUpdateInfo oldEntry,
    input logic `VADDR_BUS pc,
    input FsqIdxInfo fsqInfo,
    input logic `N(`PREDICTION_WIDTH) normalOffset,
    input BranchType br_type,
    input logic pred_error,
    input logic exception,
`ifdef RVC
    input logic rvc,
    input logic `N(`SLOT_NUM) slot_rvc, // 分支槽的前一条指令是否为rvc
    input logic rd_rvc, // 分支预测错误的前一条指令是否为rvc
`endif
    input logic `VADDR_BUS target,
    input logic `N(`SLOT_NUM) predTaken,
    input logic taken,
    output BTBUpdateInfo updateEntry,
    output logic `N(`SLOT_NUM) allocSlot,
    output logic `N(`SLOT_NUM) realTaken
);
    // 如果不是分支指令，那么插入tailSlot
    // 如果是分支指令,判断是否有空位
    // 如果有空位则在空位中插入
    // 否则将比他大的指令踢出去
    // 踢出去的规则：
    // 1. 当包含两条分支指令时，第三条指令插入时判断三者大小关系
    //   假设存在两条指令A,B,要插入的指令为I
    //   如果当前为I, A, B,那么将I插入B中，并且此时fthAddr为B
    //   如果BIA,那么将I插入A，fthAddr为A
    //   如果为ABI,那么不插入，并且fthAddr为I

    logic `N(`SLOT_NUM) free, free_p, oldest, equal, we;
    logic `ARRAY(`SLOT_NUM+1, `PREDICTION_WIDTH) offsets;
    logic `N(`PREDICTION_WIDTH) oldestOffset;
    logic `N(`SLOT_NUM+1) oldestDecode;
    logic `N(`SLOT_NUM) taken_ext;
    logic `N(`SLOT_NUM) entry_ens;
    logic `N(`SLOT_NUM) predAlloc, predOldAlloc, slotAlloc;
    logic `ARRAY(`SLOT_NUM, `SLOT_NUM) slotOldAlloc;
    logic `N(`SLOT_NUM) allocOldest;
generate
    for(genvar i=0; i<`SLOT_NUM-1; i++)begin
        assign free[i] = !entry_ens[i];
        assign offsets[i] = oldEntry.slots[i].offset;
        assign equal[i] = entry_ens[i] && oldEntry.slots[i].offset == fsqInfo.offset;
        assign entry_ens[i] = oldEntry.slots[i].en;
    end
endgenerate
    assign we = |equal ? equal :
                |free ? free_p : oldest;
    assign taken_ext = {`SLOT_NUM{taken}};
    assign free[`SLOT_NUM-1] = !oldEntry.tailSlot.en;
    assign offsets[`SLOT_NUM-1] = oldEntry.tailSlot.offset;
    assign equal[`SLOT_NUM-1] = oldEntry.tailSlot.en && oldEntry.tailSlot.br_type == CONDITION &&  oldEntry.tailSlot.offset == fsqInfo.offset;
    assign offsets[`SLOT_NUM] = fsqInfo.offset;
    assign entry_ens[`SLOT_NUM-1] = oldEntry.tailSlot.en;
    PRSelector #(`SLOT_NUM) selector_free (free, free_p);

    typedef struct packed {
        logic `N($clog2(`SLOT_NUM)+1) idx;
`ifdef RVC
        logic rvc;
`endif
    } OldestInfo;
    OldestInfo `N(`SLOT_NUM+1) selectInfos;
    OldestInfo oldestInfo;
`ifdef RVC
    for(genvar i =0; i<`SLOT_NUM; i++)begin
        assign selectInfos[i].rvc = slot_rvc[i];
    end
    assign selectInfos[`SLOT_NUM].rvc = rd_rvc;
`endif
    for(genvar i=0; i<`SLOT_NUM+1; i++)begin
        assign selectInfos[i].idx = i;
    end
    OldestSelect #(
        .RADIX(`SLOT_NUM+1),
        .WIDTH(`PREDICTION_WIDTH),
        .DATA_WIDTH($bits(OldestInfo))
    ) oldest_select (
        .cmp(offsets),
        .data_i(selectInfos),
        .cmp_o(oldestOffset),
        .data_o(oldestInfo)
    );
    Decoder #(`SLOT_NUM+1) decode_oldest(oldestInfo.idx, oldestDecode);
    assign oldest = oldestDecode[`SLOT_NUM-1: 0];

    TargetState tarState, tailTarState;
    assign tarState = target[`VADDR_SIZE-1: `JAL_OFFSET+1] > pc[`VADDR_SIZE-1: `JAL_OFFSET+1] ? TAR_OV :
                      target[`VADDR_SIZE-1: `JAL_OFFSET+1] < pc[`VADDR_SIZE-1: `JAL_OFFSET+1] ? TAR_UN : TAR_NONE;
    assign tailTarState = target[`VADDR_SIZE-1: `JALR_OFFSET+1] > pc[`VADDR_SIZE-1: `JALR_OFFSET+1] ? TAR_OV :
                      target[`VADDR_SIZE-1: `JALR_OFFSET+1] < pc[`VADDR_SIZE-1: `JALR_OFFSET+1] ? TAR_UN : TAR_NONE;
    always_comb begin
        updateEntry.en = 1'b1;
        if(br_type != CONDITION)begin
            updateEntry.slots = oldEntry.slots;
            if(&allocOldest)begin // 如果预测错误的分支是最老的则不需要更新tailSlot
                updateEntry.fthAddr = oldestOffset-{~oldestInfo.rvc, oldestInfo.rvc};
`ifdef RVC
                updateEntry.fth_rvc = oldestInfo.rvc;
`endif
                updateEntry.tailSlot = oldEntry.tailSlot;
            end
            else begin
                // updateEntry.fthAddr = fsqInfo.offset;
                updateEntry.fthAddr = `BLOCK_INST_SIZE-1;
                updateEntry.tailSlot.en = 1'b1;
                updateEntry.tailSlot.carry = ~oldEntry.tailSlot.en;
                updateEntry.tailSlot.br_type = br_type;
    `ifdef RVC
                updateEntry.tailSlot.rvc = rvc;
                updateEntry.fth_rvc = 1'b1;
    `endif
                updateEntry.tailSlot.offset = fsqInfo.offset;
                updateEntry.tailSlot.target = target[`JALR_OFFSET: 1];
                updateEntry.tailSlot.tar_state = tailTarState;
            end
        end
        else begin
            for(int i=0; i<`SLOT_NUM-1; i++)begin
                updateEntry.slots[i].en = we[i] | oldEntry.slots[i].en;
                updateEntry.slots[i].carry = (oldEntry.slots[i].carry | free_p[i]) & ~equal[i];
                updateEntry.slots[i].offset = we[i] ? fsqInfo.offset : 
                                              oldEntry.slots[i].en ? oldEntry.slots[i].offset :
                                              `BLOCK_INST_SIZE - 1;
                updateEntry.slots[i].target = we[i] & taken ? target[`JAL_OFFSET: 1] : oldEntry.slots[i].target;
                updateEntry.slots[i].tar_state = we[i] & taken ? tarState : oldEntry.slots[i].tar_state;
`ifdef RVC
                updateEntry.slots[i].rvc = we[i] ? rvc : oldEntry.slots[i].rvc;
`endif
            end
            updateEntry.tailSlot.en = we[`SLOT_NUM-1] ? 1'b1 : oldEntry.tailSlot.en;
            updateEntry.tailSlot.carry = (oldEntry.tailSlot.carry | free_p[`SLOT_NUM-1]) & ~equal[`SLOT_NUM-1];
            updateEntry.tailSlot.br_type = we[`SLOT_NUM-1] ? br_type : oldEntry.tailSlot.br_type;
            updateEntry.tailSlot.offset = we[`SLOT_NUM-1] ? fsqInfo.offset : 
                                          oldEntry.tailSlot.en ? oldEntry.tailSlot.offset :
                                          `BLOCK_INST_SIZE - 1;
            updateEntry.tailSlot.target = we[`SLOT_NUM-1] ? target[`JAL_OFFSET: 1] : oldEntry.tailSlot.target;
            updateEntry.tailSlot.tar_state = we[`SLOT_NUM-1] ? tarState : oldEntry.tailSlot.tar_state;
`ifdef RVC
            updateEntry.tailSlot.rvc = we[`SLOT_NUM-1] ? rvc : oldEntry.tailSlot.rvc;
            updateEntry.fthAddr = (~(|free)) & (~(|equal)) ? oldestOffset-{~oldestInfo.rvc, oldestInfo.rvc} : 
                                  oldEntry.en ? oldEntry.fthAddr : `BLOCK_INST_SIZE-1;
            updateEntry.fth_rvc = (~(|free)) & (~(|equal)) ? oldestInfo.rvc :
                                  oldEntry.en ? oldEntry.fth_rvc : 1'b1;
`else
            updateEntry.fthAddr = (~(|free)) & (~(|equal)) ? oldestOffset-1 : 
                                  oldEntry.en ? oldEntry.fthAddr : `BLOCK_INST_SIZE-1;
`endif
        end
    end

    always_comb begin
        if((~pred_error) | exception)begin
            realTaken = predTaken;
        end
        else if(|equal)begin
            realTaken = (equal & taken_ext);
        end
        else if(|free)begin
            realTaken = (free_p & taken_ext);
        end
        else begin
            realTaken = (oldest[`SLOT_NUM-1: 0] & taken_ext);
        end
    end

generate
    for(genvar i=0; i<`SLOT_NUM; i++)begin
        assign predAlloc[i] = ~free[i]  & (normalOffset >= offsets[i]);
        assign predOldAlloc[i] = ~free[i] & ((fsqInfo.offset > offsets[i]) | equal[i]);
        assign allocOldest[i] = ~free[i] & (fsqInfo.offset > offsets[i]);
        for(genvar j=0; j<`SLOT_NUM; j++)begin
            if(i == j)begin
                assign slotOldAlloc[i][j] = equal[i];
            end
            else begin
                assign slotOldAlloc[i][j] = ~free[j] & equal[i] & (offsets[i] > offsets[j]);
            end
        end
    end
endgenerate
    ParallelOR #(`SLOT_NUM, `SLOT_NUM) or_slotOldAlloc (slotOldAlloc, slotAlloc);
    always_comb begin
        if(~pred_error | exception)begin
            allocSlot = predAlloc;
        end
        else if(|equal)begin
            allocSlot = (br_type != CONDITION) & equal[`SLOT_NUM-1] ? 
                        {1'b1, allocOldest[`SLOT_NUM-2:0] & {`SLOT_NUM-1{equal[`SLOT_NUM-1]}}} : predOldAlloc;
        end
        else if(|free)begin
            allocSlot = predOldAlloc | (br_type == CONDITION ? free_p : {1'b1, {`SLOT_NUM-1{1'b0}}});
        end
        else begin
            allocSlot = predOldAlloc | (br_type == CONDITION ? we : {1'b1, {`SLOT_NUM-1{1'b0}}});
        end
    end

endmodule