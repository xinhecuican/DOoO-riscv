VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sky130_sram_1r1w0rw_32x64_8
   CLASS BLOCK ;
   SIZE 368.26 BY 252.18 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  98.62 0.0 99.0 0.38 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  104.46 0.0 104.84 0.38 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  110.3 0.0 110.68 0.38 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  116.14 0.0 116.52 0.38 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  121.98 0.0 122.36 0.38 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  127.82 0.0 128.2 0.38 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  133.66 0.0 134.04 0.38 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  139.5 0.0 139.88 0.38 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  145.34 0.0 145.72 0.38 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  151.18 0.0 151.56 0.38 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  157.02 0.0 157.4 0.38 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  162.86 0.0 163.24 0.38 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  168.7 0.0 169.08 0.38 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  174.54 0.0 174.92 0.38 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  180.38 0.0 180.76 0.38 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  186.22 0.0 186.6 0.38 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  192.06 0.0 192.44 0.38 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  197.9 0.0 198.28 0.38 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  203.74 0.0 204.12 0.38 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  209.58 0.0 209.96 0.38 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  215.42 0.0 215.8 0.38 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  221.26 0.0 221.64 0.38 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  227.1 0.0 227.48 0.38 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  232.94 0.0 233.32 0.38 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  238.78 0.0 239.16 0.38 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  244.62 0.0 245.0 0.38 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  250.46 0.0 250.84 0.38 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  256.3 0.0 256.68 0.38 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  262.14 0.0 262.52 0.38 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  267.98 0.0 268.36 0.38 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  273.82 0.0 274.2 0.38 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  279.66 0.0 280.04 0.38 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 107.58 0.38 107.96 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 116.08 0.38 116.46 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 121.72 0.38 122.1 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 130.22 0.38 130.6 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 136.275 0.38 136.655 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 144.675 0.38 145.055 ;
      END
   END addr0[5]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  306.53 0.0 306.91 0.38 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  302.175 0.0 302.555 0.38 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  305.84 0.0 306.22 0.38 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  302.865 0.0 303.245 0.38 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  303.555 0.0 303.935 0.38 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  304.3 0.0 304.68 0.38 ;
      END
   END addr1[5]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 14.87 0.38 15.25 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  367.88 237.075 368.26 237.455 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  30.26 0.0 30.64 0.38 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  337.62 251.8 338.0 252.18 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  75.26 0.0 75.64 0.38 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  81.1 0.0 81.48 0.38 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  86.94 0.0 87.32 0.38 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  92.78 0.0 93.16 0.38 ;
      END
   END wmask0[3]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  134.445 251.8 134.825 252.18 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  139.415 251.8 139.795 252.18 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  140.685 251.8 141.065 252.18 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  145.655 251.8 146.035 252.18 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  146.925 251.8 147.305 252.18 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  151.895 251.8 152.275 252.18 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  153.165 251.8 153.545 252.18 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  158.135 251.8 158.515 252.18 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  159.405 251.8 159.785 252.18 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  164.375 251.8 164.755 252.18 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  165.645 251.8 166.025 252.18 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  170.615 251.8 170.995 252.18 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  171.885 251.8 172.265 252.18 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  176.855 251.8 177.235 252.18 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  178.125 251.8 178.505 252.18 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  183.095 251.8 183.475 252.18 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  184.365 251.8 184.745 252.18 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  189.335 251.8 189.715 252.18 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  190.605 251.8 190.985 252.18 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  195.575 251.8 195.955 252.18 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  196.845 251.8 197.225 252.18 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  201.815 251.8 202.195 252.18 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  203.085 251.8 203.465 252.18 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  208.055 251.8 208.435 252.18 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  209.325 251.8 209.705 252.18 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  214.295 251.8 214.675 252.18 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  215.565 251.8 215.945 252.18 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  220.535 251.8 220.915 252.18 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  221.805 251.8 222.185 252.18 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  226.775 251.8 227.155 252.18 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  228.045 251.8 228.425 252.18 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  233.015 251.8 233.395 252.18 ;
      END
   END dout1[31]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  0.0 250.44 368.26 252.18 ;
         LAYER met3 ;
         RECT  0.0 0.0 368.26 1.74 ;
         LAYER met4 ;
         RECT  366.52 0.0 368.26 252.18 ;
         LAYER met4 ;
         RECT  0.0 0.0 1.74 252.18 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  3.48 3.48 5.22 248.7 ;
         LAYER met3 ;
         RECT  3.48 3.48 364.78 5.22 ;
         LAYER met4 ;
         RECT  363.04 3.48 364.78 248.7 ;
         LAYER met3 ;
         RECT  3.48 246.96 364.78 248.7 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 367.64 251.56 ;
   LAYER  met2 ;
      RECT  0.62 0.62 367.64 251.56 ;
   LAYER  met3 ;
      RECT  0.98 106.98 367.64 108.56 ;
      RECT  0.62 108.56 0.98 115.48 ;
      RECT  0.62 117.06 0.98 121.12 ;
      RECT  0.62 122.7 0.98 129.62 ;
      RECT  0.62 131.2 0.98 135.675 ;
      RECT  0.62 137.255 0.98 144.075 ;
      RECT  0.62 15.85 0.98 106.98 ;
      RECT  0.98 108.56 367.28 236.475 ;
      RECT  0.98 236.475 367.28 238.055 ;
      RECT  367.28 108.56 367.64 236.475 ;
      RECT  0.62 145.655 0.98 249.84 ;
      RECT  367.28 238.055 367.64 249.84 ;
      RECT  0.62 2.34 0.98 14.27 ;
      RECT  0.98 2.34 2.88 2.88 ;
      RECT  0.98 2.88 2.88 5.82 ;
      RECT  0.98 5.82 2.88 106.98 ;
      RECT  2.88 2.34 365.38 2.88 ;
      RECT  2.88 5.82 365.38 106.98 ;
      RECT  365.38 2.34 367.64 2.88 ;
      RECT  365.38 2.88 367.64 5.82 ;
      RECT  365.38 5.82 367.64 106.98 ;
      RECT  0.98 238.055 2.88 246.36 ;
      RECT  0.98 246.36 2.88 249.3 ;
      RECT  0.98 249.3 2.88 249.84 ;
      RECT  2.88 238.055 365.38 246.36 ;
      RECT  2.88 249.3 365.38 249.84 ;
      RECT  365.38 238.055 367.28 246.36 ;
      RECT  365.38 246.36 367.28 249.3 ;
      RECT  365.38 249.3 367.28 249.84 ;
   LAYER  met4 ;
      RECT  98.02 0.98 99.6 251.56 ;
      RECT  99.6 0.62 103.86 0.98 ;
      RECT  105.44 0.62 109.7 0.98 ;
      RECT  111.28 0.62 115.54 0.98 ;
      RECT  117.12 0.62 121.38 0.98 ;
      RECT  122.96 0.62 127.22 0.98 ;
      RECT  128.8 0.62 133.06 0.98 ;
      RECT  134.64 0.62 138.9 0.98 ;
      RECT  140.48 0.62 144.74 0.98 ;
      RECT  146.32 0.62 150.58 0.98 ;
      RECT  152.16 0.62 156.42 0.98 ;
      RECT  158.0 0.62 162.26 0.98 ;
      RECT  163.84 0.62 168.1 0.98 ;
      RECT  169.68 0.62 173.94 0.98 ;
      RECT  175.52 0.62 179.78 0.98 ;
      RECT  181.36 0.62 185.62 0.98 ;
      RECT  187.2 0.62 191.46 0.98 ;
      RECT  193.04 0.62 197.3 0.98 ;
      RECT  198.88 0.62 203.14 0.98 ;
      RECT  204.72 0.62 208.98 0.98 ;
      RECT  210.56 0.62 214.82 0.98 ;
      RECT  216.4 0.62 220.66 0.98 ;
      RECT  222.24 0.62 226.5 0.98 ;
      RECT  228.08 0.62 232.34 0.98 ;
      RECT  233.92 0.62 238.18 0.98 ;
      RECT  239.76 0.62 244.02 0.98 ;
      RECT  245.6 0.62 249.86 0.98 ;
      RECT  251.44 0.62 255.7 0.98 ;
      RECT  257.28 0.62 261.54 0.98 ;
      RECT  263.12 0.62 267.38 0.98 ;
      RECT  268.96 0.62 273.22 0.98 ;
      RECT  274.8 0.62 279.06 0.98 ;
      RECT  280.64 0.62 301.575 0.98 ;
      RECT  99.6 0.98 337.02 251.2 ;
      RECT  337.02 0.98 338.6 251.2 ;
      RECT  31.24 0.62 74.66 0.98 ;
      RECT  76.24 0.62 80.5 0.98 ;
      RECT  82.08 0.62 86.34 0.98 ;
      RECT  87.92 0.62 92.18 0.98 ;
      RECT  93.76 0.62 98.02 0.98 ;
      RECT  99.6 251.2 133.845 251.56 ;
      RECT  135.425 251.2 138.815 251.56 ;
      RECT  141.665 251.2 145.055 251.56 ;
      RECT  147.905 251.2 151.295 251.56 ;
      RECT  154.145 251.2 157.535 251.56 ;
      RECT  160.385 251.2 163.775 251.56 ;
      RECT  166.625 251.2 170.015 251.56 ;
      RECT  172.865 251.2 176.255 251.56 ;
      RECT  179.105 251.2 182.495 251.56 ;
      RECT  185.345 251.2 188.735 251.56 ;
      RECT  191.585 251.2 194.975 251.56 ;
      RECT  197.825 251.2 201.215 251.56 ;
      RECT  204.065 251.2 207.455 251.56 ;
      RECT  210.305 251.2 213.695 251.56 ;
      RECT  216.545 251.2 219.935 251.56 ;
      RECT  222.785 251.2 226.175 251.56 ;
      RECT  229.025 251.2 232.415 251.56 ;
      RECT  233.995 251.2 337.02 251.56 ;
      RECT  307.51 0.62 365.92 0.98 ;
      RECT  338.6 251.2 365.92 251.56 ;
      RECT  2.34 0.62 29.66 0.98 ;
      RECT  2.34 0.98 2.88 2.88 ;
      RECT  2.34 2.88 2.88 249.3 ;
      RECT  2.34 249.3 2.88 251.56 ;
      RECT  2.88 0.98 5.82 2.88 ;
      RECT  2.88 249.3 5.82 251.56 ;
      RECT  5.82 0.98 98.02 2.88 ;
      RECT  5.82 2.88 98.02 249.3 ;
      RECT  5.82 249.3 98.02 251.56 ;
      RECT  338.6 0.98 362.44 2.88 ;
      RECT  338.6 2.88 362.44 249.3 ;
      RECT  338.6 249.3 362.44 251.2 ;
      RECT  362.44 0.98 365.38 2.88 ;
      RECT  362.44 249.3 365.38 251.2 ;
      RECT  365.38 0.98 365.92 2.88 ;
      RECT  365.38 2.88 365.92 249.3 ;
      RECT  365.38 249.3 365.92 251.2 ;
   END
END    sky130_sram_1r1w0rw_32x64_8
END    LIBRARY
