`ifndef ARCH_H
`define ARCH_H

`define RV32I
`define ZICSR
`define DIFFTEST
`endif
