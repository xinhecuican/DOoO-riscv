`include "../../defines/defines.svh"

// btb update: idx, updateEntry
// tage update: pred, pred error

module FSQ (
    input logic clk,
    input logic rst,
    BpuFsqIO.fsq bpu_fsq_io,
    FsqCacheIO.fsq fsq_cache_io,
    PreDecodeRedirect.redirect pd_redirect,
    FsqBackendIO.fsq fsq_back_io,
    CommitBus commitBus,
    FrontendCtrl frontendCtrl
);
    logic `N(`FSQ_WIDTH) search_head, commit_head, tail, write_index, tail_n1, n_commit_head;
    logic `N(`FSQ_WIDTH) write_tail;
    logic `N(`FSQ_WIDTH) squashIdx;
    logic full, enqueue, dequeue;
    logic queue_we;
    logic last_search;
    logic empty;
    logic cache_req_ok;
    BTBEntry oldEntry, updateEntry;
    logic `N(`BLOCK_INST_SIZE) predErrorVec `N(`FSQ_SIZE);
    logic directionTable `N(`FSQ_SIZE);
    logic direction, hdir;
    FetchStream commitStream;
    logic `ARRAY(2, `BLOCK_INST_SIZE) commitVec, streamVec;
    logic `ARRAY(`COMMIT_WIDTH, `BLOCK_INST_SIZE * 2) commitOffsetExpand;
    logic commitValid;
    BTBEntry commitUpdateEntry;
    

    assign tail_n1 = tail + 1;
    assign write_tail = bpu_fsq_io.redirect ? bpu_fsq_io.stream_idx : tail;
    assign queue_we = bpu_fsq_io.en;
    assign write_index = bpu_fsq_io.redirect ? bpu_fsq_io.stream_idx : tail;
    MPRAM #(
        .WIDTH($bits(FetchStream)),
        .DEPTH(`FSQ_SIZE),
        .READ_PORT(1+`ALU_SIZE + 1),
        .WRITE_PORT(1)
    ) fs_queue(
        .clk(clk),
        .en({(1+`ALU_SIZE+1){1'b1}}),
        .we(queue_we),
        .waddr(write_tail),
        .raddr({search_head, fsq_back_io.fsqIdx, n_commit_head}),
        .wdata(bpu_fsq_io.prediction.stream),
        .rdata({fsq_cache_io.stream, fsq_back_io.streams, commitStream})
    );

    RedirectInfo redirect_regs `N(`FSQ_SIZE);
    RedirectInfo u_redirectInfo, c_redirectInfo;


    assign squashIdx = fsq_back_io.redirect.en ? fsq_back_io.redirect.fsqInfo.idx : pd_redirect.fsqIdx;
    assign u_redirectInfo = redirect_regs[squashIdx];
    always_ff @(posedge clk)begin
        if(queue_we)begin
            redirect_regs[write_tail] <= bpu_fsq_io.prediction.redirect_info;
        end
    end

    MPRAM #(
        .WIDTH($bits(BTBEntry)),
        .DEPTH(`FSQ_SIZE),
        .READ_PORT(1),
        .WRITE_PORT(1)
    ) btb_ram (
        .clk(clk),
        .en(1'b1),
        .raddr(n_commit_head),
        .rdata(oldEntry),
        .we(queue_we),
        .waddr(write_tail),
        .wdata(bpu_fsq_io.prediction.btbEntry)
    );

    PredictionMeta updateMeta;
    MPRAM #(
        .WIDTH($bits(PredictionMeta)),
        .DEPTH(`FSQ_SIZE),
        .READ_PORT(1),
        .WRITE_PORT(1)
    ) meta_ram (
        .clk(clk),
        .en(1'b1),
        .raddr(commit_head),
        .rdata(updateMeta),
        .we(bpu_fsq_io.lastStage),
        .waddr(bpu_fsq_io.lastStageIdx),
        .wdata(bpu_fsq_io.lastStageMeta)
    );

    typedef struct packed {
        logic `N(2) condNum;
        logic `N(`SLOT_NUM) condHist;
        logic `N(`SLOT_NUM) condValid;
        logic `ARRAY(`SLOT_NUM, `PREDICTION_WIDTH) offsets;
    } PredictionInfo;

    PredictionInfo predictionInfos `N(`FSQ_SIZE);
    PredictionInfo pd_wr_info;
    logic `N(2) condNum;
    logic `N(`SLOT_NUM) condSmallNum;
    logic `N(`SLOT_NUM) condSmallNumAll;
    logic redirectIsCond;
    PredictionInfo redirectPredInfo;
    PredictionInfo pd_predInfo;
    PredictionInfo u_predInfo;

    assign pd_wr_info.condNum = bpu_fsq_io.prediction.cond_num;
    assign pd_wr_info.condHist = bpu_fsq_io.prediction.predTaken;
    BTBEntry predEntry;
    assign predEntry = bpu_fsq_io.prediction.btbEntry;
generate
    for(genvar i=0; i<`SLOT_NUM-1; i++)begin
        assign pd_wr_info.offsets[i] = predEntry.slots[i].offset;
    end
    assign pd_wr_info.condValid = bpu_fsq_io.prediction.cond_valid;
    assign pd_wr_info.offsets[`SLOT_NUM-1] = predEntry.tailSlot.offset;
endgenerate

    always_ff @(posedge clk)begin
        if(rst == `RST)begin
            predictionInfos <= '{default: 0};
        end
        else begin
            if(queue_we)begin
                predictionInfos[write_tail] <= pd_wr_info;
            end
        end
    end

    assign fsq_cache_io.en = search_head != tail || full;
    assign fsq_cache_io.abandon = bpu_fsq_io.redirect;
    assign fsq_cache_io.abandonIdx = bpu_fsq_io.prediction.stream_idx;
    assign fsq_cache_io.flush = pd_redirect.en | fsq_back_io.redirect.en;
    assign fsq_cache_io.stall = frontendCtrl.ibuf_full;
    assign bpu_fsq_io.stream_idx = tail;
    assign bpu_fsq_io.stream_dir = direction;
    assign bpu_fsq_io.stall = full;
    assign cache_req_ok = fsq_cache_io.en & fsq_cache_io.ready;

    // logic `N(`SLOT_NUM) condFree;
    // PEncoder #(`SLOT_NUM) encoder_condFree({~oldEntry.slots[0].en, ~oldEntry.tailSlot.en}, condFree);

    assign enqueue = bpu_fsq_io.en;
    assign dequeue = pd_redirect.en | cache_req_ok | (bpu_fsq_io.redirect && (tail != bpu_fsq_io.stream_idx));

    CondPredInfo redirectCondInfo, pd_condInfo;
    assign pd_predInfo = predictionInfos[pd_redirect.fsqIdx];
    assign redirectPredInfo = predictionInfos[fsq_back_io.redirect.fsqInfo.idx];

    assign pd_condInfo.condNum = pd_predInfo.condNum;
    assign pd_condInfo.taken = |(pd_predInfo.condValid & pd_predInfo.condHist);
generate
    for(genvar i=0; i<`SLOT_NUM; i++)begin
        assign condSmallNum[i] = redirectPredInfo.condValid[i] & (redirectPredInfo.offsets[i] < fsq_back_io.redirect.fsqInfo.offset);
    end
endgenerate
    assign redirectIsCond = fsq_back_io.redirect.en & fsq_back_io.redirect.br_type == CONDITION;
    assign condSmallNumAll = condSmallNum[0] + condSmallNum[1];
    always_comb begin
        if(redirectIsCond)begin
            if(condSmallNumAll < `SLOT_NUM)begin
                redirectCondInfo.condNum = condSmallNumAll + 1;
                redirectCondInfo.taken = fsq_back_io.redirect.taken;
            end
            else begin
                redirectCondInfo.condNum = `SLOT_NUM;
                redirectCondInfo.taken = 0;
            end
        end
        else begin
            redirectCondInfo.condNum = condSmallNumAll;
            redirectCondInfo.taken = 0;
        end
    end

    assign n_commit_head = commitValid ? commit_head + 1 : commit_head;
    assign full = commit_head == tail && (hdir ^ direction);
    always_ff @(posedge clk)begin
        last_search <= search_head == tail && fsq_cache_io.en;
        bpu_fsq_io.squash <= pd_redirect.en | fsq_back_io.redirect.en;
        bpu_fsq_io.squashInfo.redirectInfo <= u_redirectInfo;
        bpu_fsq_io.squashInfo.target_pc <= fsq_back_io.redirect.en ? fsq_back_io.redirect.target : pd_redirect.redirect_addr;
        bpu_fsq_io.squashInfo.predInfo <= fsq_back_io.redirect.en ? redirectPredInfo : pd_predInfo;
        bpu_fsq_io.squashInfo.br_type <= fsq_back_io.redirect.en ? fsq_back_io.redirect.br_type : DIRECT;
        bpu_fsq_io.squashInfo.ras_type <= fsq_back_io.redirect.en ? fsq_back_io.redirect.ras_type : NONE;
        if(rst == `RST)begin
            search_head <= 0;
            commit_head <= 0;
            tail <= 0;
            predErrorVec <= '{default: 0};
        end
        else begin
            if(fsq_back_io.redirect.en)begin
                search_head <= fsq_back_io.redirect.fsqInfo.idx;
            end
            else if(!frontendCtrl.ibuf_full) begin
                if(pd_redirect.en)begin
                    search_head <= pd_redirect.fsqIdx;
                end
                else if(cache_req_ok)begin
                    search_head <= search_head + 1;
                end
            end

            if(fsq_back_io.redirect.en)begin
                tail <= fsq_back_io.redirect.fsqInfo.idx;
            end
            else if(pd_redirect.en)begin
                tail <= pd_redirect.fsqIdx;
            end
            else if(bpu_fsq_io.redirect)begin
                tail <= bpu_fsq_io.stream_idx + 1;
            end
            else if(bpu_fsq_io.en)begin
                tail <= tail_n1;
            end

            commit_head <= n_commit_head;

            if(fsq_back_io.redirect.en)begin
                predErrorVec[fsq_back_io.redirect.fsqInfo.idx] <= predErrorVec[fsq_back_io.redirect.fsqInfo.idx] | (1 << fsq_back_io.redirect.fsqInfo.offset);
            end
        end
    end

    logic `N(`FSQ_WIDTH) redirect_dir_idx;
    assign redirect_dir_idx = fsq_back_io.redirect.en ? fsq_back_io.redirect.fsqInfo.idx : pd_redirect.fsqIdx;
    always_ff @(posedge clk)begin
        for(int i=0; i<`ALU_SIZE; i++)begin
            fsq_back_io.directions[i] <= directionTable[fsq_back_io.fsqIdx[i]];
        end

        if(rst == `RST)begin
            direction <= 0;
            hdir <= 0;
            directionTable <= '{default: 0};
        end
        else begin
            if(pd_redirect.en | fsq_back_io.redirect.en)begin
                direction <= directionTable[redirect_dir_idx];
            end
            else if(bpu_fsq_io.redirect)begin
                direction <= bpu_fsq_io.stream_dir;
            end
            else if(bpu_fsq_io.en)begin
                direction <= tail[`FSQ_WIDTH-1] ^ tail_n1[`FSQ_WIDTH-1] ? ~direction : direction;
            end
            if(commitValid)begin
                hdir <= commit_head[`FSQ_WIDTH-1] ^ n_commit_head[`FSQ_WIDTH-1] ? ~hdir : hdir;
            end

            if(bpu_fsq_io.en)begin
                directionTable[tail] <= direction;
            end
        end
    end

    typedef struct packed {
        logic en;
        logic taken;
        BranchType br_type;
        RasType ras_type;
        logic `N(`VADDR_SIZE) target;
        logic `N(`PREDICTION_WIDTH) offset;
    } WBInfo;

    WBInfo wbInfos `N(`RAS_SIZE);
    BackendRedirectInfo rd;
    assign rd = fsq_back_io.redirect;
    always_ff @(posedge clk)begin
        if(rst == `RST)begin
            wbInfos <= '{default: 0};
        end
        else begin
            if(rd.en)begin
                wbInfos[rd.fsqInfo.idx] <= {1'b1, rd.taken, rd.br_type, rd.ras_type, rd.target, rd.fsqInfo.offset};
            end
        end
    end

    assign streamVec = (1 << (commitStream.size + 1)) - 1;
    assign commitValid = ((streamVec & commitVec[tail[0]]) == streamVec) |
                         ((streamVec & predErrorVec[tail]) != 0);
generate
    for(genvar i=0; i<`COMMIT_WIDTH; i++)begin
        logic `N(`BLOCK_INST_SIZE) commitOffsetDecode;
        Decoder #(`BLOCK_INST_SIZE) decoder_commit_offset (commitBus.fsqInfo[i].offset, commitOffsetDecode);
        assign commitOffsetExpand[i] =  {{`BLOCK_INST_SIZE{commitBus.fsqInfo[i].idx[0] & commitBus.en[i]}} & commitOffsetDecode,
                                        {`BLOCK_INST_SIZE{~commitBus.fsqInfo[i].idx[0] & commitBus.en[i]}} & commitOffsetDecode};
    end
endgenerate

    always_ff @(posedge clk)begin
        if(rst == `RST)begin
            commitVec <= 0;
        end
        else begin
            commitVec <= (commitVec | (|commitOffsetExpand));
        end
    end
    FsqIdxInfo commitFsqInfo;
    logic `N(`SLOT_NUM) realTaken, allocSlot;
    assign u_predInfo = predictionInfos[commitFsqInfo.idx];
    assign commitFsqInfo.idx = tail;
    assign commitFsqInfo.offset = wbInfos[tail].offset;
    BTBEntryGen commit_btb_entry_gen (
        .oldEntry(oldEntry),
        .pc(commitStream.start_addr),
        .fsqInfo(commitFsqInfo),
        .br_type(wbInfos[tail].br_type),
        .ras_type(wbInfos[tail].ras_type),
        .target(wbInfos[tail].target),
        .taken(wbInfos[tail].taken),
        .predTaken(u_predInfo.condHist),
        .updateEntry(commitUpdateEntry),
        .realTaken(realTaken),
        .allocSlot(allocSlot)
    );

    BranchUpdateInfo updateInfo;
    assign updateInfo.start_addr = commitStream.start_addr;
    assign updateInfo.target_pc = wbInfos[tail].target;
    assign updateInfo.redirectInfo = c_redirectInfo;
    assign updateInfo.btbEntry = commitUpdateEntry;
    assign updateInfo.meta = updateMeta;
    assign updateInfo.realTaken = realTaken;
    assign updateInfo.allocSlot = allocSlot;
    always_ff @(posedge clk)begin
        bpu_fsq_io.update <= commitValid;
        bpu_fsq_io.updateInfo <= updateInfo;
    end
endmodule

module BTBEntryGen(
    input BTBEntry oldEntry,
    input logic `VADDR_BUS pc,
    input FsqIdxInfo fsqInfo,
    input BranchType br_type,
    input RasType ras_type,
    input logic `VADDR_BUS target,
    input logic `N(`SLOT_NUM) predTaken,
    input logic taken,
    output BTBEntry updateEntry,
    output logic `N(`SLOT_NUM) allocSlot,
    output logic `N(`SLOT_NUM) realTaken
);
    // 如果不是分支指令，那么插入tailSlot
    // 如果是分支指令,判断是否有空位
    // 如果有空位则在空位中插入
    // 否则将比他大的指令踢出去
    // 踢出去的规则：
    // 1. 当包含两条分支指令时，第三条指令插入时判断三者大小关系
    //   假设存在两条指令A,B,要插入的指令为I
    //   如果当前为I, A, B,那么将I插入B中，并且此时fthAddr为B
    //   如果BIA,那么将I插入A，fthAddr为A
    //   如果为ABI,那么不插入，并且fthAddr为I

    logic `N(`SLOT_NUM) free, free_p, oldest, equal, we;
    logic `ARRAY(`SLOT_NUM+1, `PREDICTION_WIDTH) offsets;
    logic `ARRAY(`SLOT_NUM+1, $clog2(`SLOT_NUM+1)) idx;
    logic `N(`PREDICTION_WIDTH) oldestOffset;
    logic `N($clog2(`SLOT_NUM+1)) oldestIdx;
    logic `N(`SLOT_NUM+1) oldestDecode;
    logic `N(`SLOT_NUM) taken_ext;
generate
    for(genvar i=0; i<`SLOT_NUM-1; i++)begin
        assign free[i] = !oldEntry.slots[i].en;
        assign offsets[i] = oldEntry.slots[i].offset;
        assign equal[i] = oldEntry.slots[i].en && oldEntry.slots[i].offset == fsqInfo.offset;
    end
endgenerate
    assign we = |equal ? equal :
                |free ? free_p : oldest;
    assign taken_ext = {`SLOT_NUM{taken}};
    assign realTaken = |equal ? (equal & taken_ext) | (~equal & predTaken) :
                       |free ? (free & taken_ext) | (~free & predTaken) :
                       (oldest[`SLOT_NUM-1: 0] & taken_ext) | (~oldest[`SLOT_NUM-1: 0] & predTaken);
    assign allocSlot = ~(|free) & ~(|equal) & br_type == CONDITION ? oldest : 0;
    assign free[`SLOT_NUM-1] = !oldEntry.tailSlot.en;
    assign offsets[`SLOT_NUM-1] = oldEntry.tailSlot.offset;
    assign equal[`SLOT_NUM-1] = oldEntry.tailSlot.en && oldEntry.tailSlot.br_type == CONDITION &&  oldEntry.tailSlot.offset == fsqInfo.offset;
    assign offsets[`SLOT_NUM] = fsqInfo.offset;
    PSelector #(`SLOT_NUM) selector_free (free, free_p);
    for(genvar i=0; i<`SLOT_NUM+1; i++)begin
        assign idx[i] = i;
    end
    OldestSelect #(
        .RADIX(`SLOT_NUM+1),
        .WIDTH(`PREDICTION_WIDTH),
        .DATA_WIDTH($clog2(`SLOT_NUM+1))
    ) oldest_select (
        .cmp(offsets),
        .data_i(idx),
        .cmp_o(oldestOffset),
        .data_o(oldestIdx)
    );
    Decoder #(`SLOT_NUM+1) decode_oldest(oldestIdx, oldestDecode);
    assign oldest = oldestDecode[`SLOT_NUM-1: 0];


    always_comb begin
        if(br_type != CONDITION)begin
            updateEntry.en = 1'b1;
            updateEntry.tag = pc`BTB_TAG_BUS;
            updateEntry.fthAddr = fsqInfo.offset;

            updateEntry.slots = oldEntry.slots;
            updateEntry.tailSlot.en = 1'b1;
            updateEntry.tailSlot.carry = ~oldEntry.tailSlot.en;
            updateEntry.tailSlot.br_type = br_type;
            updateEntry.tailSlot.ras_type = ras_type;
            updateEntry.tailSlot.offset = fsqInfo.offset;
            updateEntry.tailSlot.target = target;
        end
        else begin
            for(int i=0; i<`SLOT_NUM-1; i++)begin
                updateEntry.slots[i].en = we[i] | oldEntry.slots[i].en;
                updateEntry.slots[i].carry = (updateEntry.slots[i].carry | free_p[i]) & ~equal[i];
                updateEntry.slots[i].offset = we[i] ? offsets[i] : oldEntry.slots[i].offset;
                updateEntry.slots[i].target = we[i] ? target : oldEntry.slots[i].target;
            end
            updateEntry.tailSlot.en = we[`SLOT_NUM-1] ? 1'b1 : oldEntry.tailSlot.en;
            updateEntry.tailSlot.carry = (updateEntry.tailSlot.carry | free_p[`SLOT_NUM-1]) & ~equal[`SLOT_NUM-1];
            updateEntry.tailSlot.br_type = we[`SLOT_NUM-1] ? br_type : oldEntry.tailSlot.br_type;
            updateEntry.tailSlot.ras_type = we[`SLOT_NUM-1] ? ras_type : oldEntry.tailSlot.ras_type;
            updateEntry.tailSlot.offset = we[`SLOT_NUM-1] ? offsets[`SLOT_NUM-1] : oldEntry.tailSlot.offset;
            updateEntry.tailSlot.target = we[`SLOT_NUM-1] ? target : oldEntry.tailSlot.target;

            updateEntry.en = 1'b1;
            updateEntry.tag = pc`BTB_TAG_BUS;
            updateEntry.fthAddr = (~(|free)) & (~(|equal)) ? oldestOffset-1 : oldEntry.fthAddr;
        end
    end


endmodule