`ifndef ARCH_H
`define ARCH_H

`define RV32I
`define DIFFTEST

`define EXT_M
`include "predefine.svh"
// `ifdef ZICSR
// parameter HAS_ZICSR=1;
// `else
// parameter HAS_ZICSR=0;
// `endif
`endif
