`ifndef ARCH_H
`define ARCH_H

`define RV32I
`define DIFFTEST
`endif
