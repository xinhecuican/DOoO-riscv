`ifndef ARCH_H
`define ARCH_H

`define RV32I
`define RVM
`define RVA
`define RVF
`define RVC
`define DIFFTEST

`define EXT_FENCEI

`define FEAT_LINKRAS
`define FEAT_SC
`define FEAT_ITTAGE_REGION

// `define SYNTH_VIVADO

`include "predefine.svh"
`endif
