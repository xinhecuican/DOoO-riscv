`ifndef DEFINES_SVH
`define DEFINES_SVH
`include "interfaces.svh"
`include "functions.svh"
`include "debug.svh"
`include "postdefine.svh"
`endif
