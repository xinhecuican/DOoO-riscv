`ifndef DEFINES_SVH
`define DEFINES_SVH
`include "interfaces.svh"

`endif