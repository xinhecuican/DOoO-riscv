`ifndef REG_SVH
`define REG_SVH

`define x0 5'h0
`define ra 5'h1
`define sp 5'h2
`define gp 5'h3
`define tp 5'h4
`define t0 5'h5
`define t1 5'h6
`define t2 5'h7
`define s0 5'h8
`define fp 5'h8
`define s1 5'h9
`define a0 5'ha
`define a1 5'hb
`define a2 5'hc
`define a3 5'hd
`define a4 5'he
`define a5 5'hf
`define a6 5'h10
`define a7 5'h11
`define s2 5'h12
`define s3 5'h13
`define s4 5'h14
`define s5 5'h15
`define s6 5'h16
`define s7 5'h17
`define s8 5'h18
`define s9 5'h19
`define a10 5'h1a
`define a11 5'h1b
`define t3 5'h1c
`define t4 5'h1d
`define t5 5'h1e
`define t6 5'h1f

`endif