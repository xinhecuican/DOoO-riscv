`include "../../defines/defines.svh"

module IFU (
    input logic clk,
    input logic rst,
    ICacheAxi.cache axi_io,
    IfuBackendIO.ifu ifu_backend_io,
    FsqBackendIO.backend fsq_back_io,
    CommitBus commitBus
);
    BpuFsqIO bpu_fsq_io;
    FsqCacheIO fsq_cache_io;
    CachePreDecodeIO cache_pd_io;
    PreDecodeRedirect pd_redirect;
    PreDecodeIBufferIO pd_ibuffer_io;
    FetchBundle fetchBundle;
    FrontendCtrl frontendCtrl;

    assign ifu_backend_io.fetchBundle = fetchBundle;
    assign frontendCtrl.redirect = fsq_back_io.redirect.en;
    BranchPredictor branch_predictor(.*);
    FSQ fsq(.*);
    ICache icache(.*);
    PreDecode predecode(.*);
    InstBuffer instBuffer(.*,
                          .full(frontendCtrl.ibuf_full));
endmodule
