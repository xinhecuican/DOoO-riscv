VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sky130_sram_1r1w0rw_68x256
   CLASS BLOCK ;
   SIZE 777.18 BY 383.405 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  113.94 0.0 114.32 0.38 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  119.78 0.0 120.16 0.38 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  125.62 0.0 126.0 0.38 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  131.46 0.0 131.84 0.38 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  137.3 0.0 137.68 0.38 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  143.14 0.0 143.52 0.38 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  148.98 0.0 149.36 0.38 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  154.82 0.0 155.2 0.38 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  160.66 0.0 161.04 0.38 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  166.5 0.0 166.88 0.38 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  172.34 0.0 172.72 0.38 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  178.18 0.0 178.56 0.38 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  184.02 0.0 184.4 0.38 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  189.86 0.0 190.24 0.38 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  195.7 0.0 196.08 0.38 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  201.54 0.0 201.92 0.38 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  207.38 0.0 207.76 0.38 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  213.22 0.0 213.6 0.38 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  219.06 0.0 219.44 0.38 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  224.9 0.0 225.28 0.38 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  230.74 0.0 231.12 0.38 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  236.58 0.0 236.96 0.38 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  242.42 0.0 242.8 0.38 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  248.26 0.0 248.64 0.38 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  254.1 0.0 254.48 0.38 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  259.94 0.0 260.32 0.38 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  265.78 0.0 266.16 0.38 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  271.62 0.0 272.0 0.38 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  277.46 0.0 277.84 0.38 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  283.3 0.0 283.68 0.38 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  289.14 0.0 289.52 0.38 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  294.98 0.0 295.36 0.38 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  300.82 0.0 301.2 0.38 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  306.66 0.0 307.04 0.38 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  312.5 0.0 312.88 0.38 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  318.34 0.0 318.72 0.38 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  324.18 0.0 324.56 0.38 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  330.02 0.0 330.4 0.38 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  335.86 0.0 336.24 0.38 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  341.7 0.0 342.08 0.38 ;
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  347.54 0.0 347.92 0.38 ;
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  353.38 0.0 353.76 0.38 ;
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  359.22 0.0 359.6 0.38 ;
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  365.06 0.0 365.44 0.38 ;
      END
   END din0[43]
   PIN din0[44]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  370.9 0.0 371.28 0.38 ;
      END
   END din0[44]
   PIN din0[45]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  376.74 0.0 377.12 0.38 ;
      END
   END din0[45]
   PIN din0[46]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  382.58 0.0 382.96 0.38 ;
      END
   END din0[46]
   PIN din0[47]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  388.42 0.0 388.8 0.38 ;
      END
   END din0[47]
   PIN din0[48]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  394.26 0.0 394.64 0.38 ;
      END
   END din0[48]
   PIN din0[49]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  400.1 0.0 400.48 0.38 ;
      END
   END din0[49]
   PIN din0[50]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  405.94 0.0 406.32 0.38 ;
      END
   END din0[50]
   PIN din0[51]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  411.78 0.0 412.16 0.38 ;
      END
   END din0[51]
   PIN din0[52]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  417.62 0.0 418.0 0.38 ;
      END
   END din0[52]
   PIN din0[53]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  423.46 0.0 423.84 0.38 ;
      END
   END din0[53]
   PIN din0[54]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  429.3 0.0 429.68 0.38 ;
      END
   END din0[54]
   PIN din0[55]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  435.14 0.0 435.52 0.38 ;
      END
   END din0[55]
   PIN din0[56]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  440.98 0.0 441.36 0.38 ;
      END
   END din0[56]
   PIN din0[57]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  446.82 0.0 447.2 0.38 ;
      END
   END din0[57]
   PIN din0[58]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  452.66 0.0 453.04 0.38 ;
      END
   END din0[58]
   PIN din0[59]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  458.5 0.0 458.88 0.38 ;
      END
   END din0[59]
   PIN din0[60]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  464.34 0.0 464.72 0.38 ;
      END
   END din0[60]
   PIN din0[61]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  470.18 0.0 470.56 0.38 ;
      END
   END din0[61]
   PIN din0[62]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  476.02 0.0 476.4 0.38 ;
      END
   END din0[62]
   PIN din0[63]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  481.86 0.0 482.24 0.38 ;
      END
   END din0[63]
   PIN din0[64]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  487.7 0.0 488.08 0.38 ;
      END
   END din0[64]
   PIN din0[65]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  493.54 0.0 493.92 0.38 ;
      END
   END din0[65]
   PIN din0[66]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  499.38 0.0 499.76 0.38 ;
      END
   END din0[66]
   PIN din0[67]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  505.22 0.0 505.6 0.38 ;
      END
   END din0[67]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  108.1 0.0 108.48 0.38 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 113.505 0.38 113.885 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 122.005 0.38 122.385 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 127.875 0.38 128.255 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 136.275 0.38 136.655 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 141.785 0.38 142.165 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 150.285 0.38 150.665 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 155.925 0.38 156.305 ;
      END
   END addr0[7]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  662.86 383.025 663.24 383.405 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  677.565 0.0 677.945 0.38 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  682.61 0.0 682.99 0.38 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  678.255 0.0 678.635 0.38 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  681.92 0.0 682.3 0.38 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  678.945 0.0 679.325 0.38 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  679.635 0.0 680.015 0.38 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  680.38 0.0 680.76 0.38 ;
      END
   END addr1[7]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 19.695 0.38 20.075 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  776.8 368.155 777.18 368.535 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  30.26 0.0 30.64 0.38 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  746.54 383.025 746.92 383.405 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  176.665 383.025 177.045 383.405 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  182.905 383.025 183.285 383.405 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  189.145 383.025 189.525 383.405 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  195.385 383.025 195.765 383.405 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  201.625 383.025 202.005 383.405 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  207.865 383.025 208.245 383.405 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  214.105 383.025 214.485 383.405 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  220.345 383.025 220.725 383.405 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  226.585 383.025 226.965 383.405 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  232.825 383.025 233.205 383.405 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  239.065 383.025 239.445 383.405 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  245.305 383.025 245.685 383.405 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  251.545 383.025 251.925 383.405 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  257.785 383.025 258.165 383.405 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  264.025 383.025 264.405 383.405 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  270.265 383.025 270.645 383.405 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  276.505 383.025 276.885 383.405 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  282.745 383.025 283.125 383.405 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  288.985 383.025 289.365 383.405 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  295.225 383.025 295.605 383.405 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  301.465 383.025 301.845 383.405 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  307.705 383.025 308.085 383.405 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  313.945 383.025 314.325 383.405 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  320.185 383.025 320.565 383.405 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  326.425 383.025 326.805 383.405 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  332.665 383.025 333.045 383.405 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  338.905 383.025 339.285 383.405 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  345.145 383.025 345.525 383.405 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  351.385 383.025 351.765 383.405 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  357.625 383.025 358.005 383.405 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  363.865 383.025 364.245 383.405 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  370.105 383.025 370.485 383.405 ;
      END
   END dout1[31]
   PIN dout1[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  376.345 383.025 376.725 383.405 ;
      END
   END dout1[32]
   PIN dout1[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  382.585 383.025 382.965 383.405 ;
      END
   END dout1[33]
   PIN dout1[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  388.825 383.025 389.205 383.405 ;
      END
   END dout1[34]
   PIN dout1[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  395.065 383.025 395.445 383.405 ;
      END
   END dout1[35]
   PIN dout1[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  401.305 383.025 401.685 383.405 ;
      END
   END dout1[36]
   PIN dout1[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  407.545 383.025 407.925 383.405 ;
      END
   END dout1[37]
   PIN dout1[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  413.785 383.025 414.165 383.405 ;
      END
   END dout1[38]
   PIN dout1[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  420.025 383.025 420.405 383.405 ;
      END
   END dout1[39]
   PIN dout1[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  426.265 383.025 426.645 383.405 ;
      END
   END dout1[40]
   PIN dout1[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  432.505 383.025 432.885 383.405 ;
      END
   END dout1[41]
   PIN dout1[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  438.745 383.025 439.125 383.405 ;
      END
   END dout1[42]
   PIN dout1[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  444.985 383.025 445.365 383.405 ;
      END
   END dout1[43]
   PIN dout1[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  451.225 383.025 451.605 383.405 ;
      END
   END dout1[44]
   PIN dout1[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  457.465 383.025 457.845 383.405 ;
      END
   END dout1[45]
   PIN dout1[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  463.705 383.025 464.085 383.405 ;
      END
   END dout1[46]
   PIN dout1[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  469.945 383.025 470.325 383.405 ;
      END
   END dout1[47]
   PIN dout1[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  476.185 383.025 476.565 383.405 ;
      END
   END dout1[48]
   PIN dout1[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  482.425 383.025 482.805 383.405 ;
      END
   END dout1[49]
   PIN dout1[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  488.665 383.025 489.045 383.405 ;
      END
   END dout1[50]
   PIN dout1[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  494.905 383.025 495.285 383.405 ;
      END
   END dout1[51]
   PIN dout1[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  501.145 383.025 501.525 383.405 ;
      END
   END dout1[52]
   PIN dout1[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  507.385 383.025 507.765 383.405 ;
      END
   END dout1[53]
   PIN dout1[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  513.625 383.025 514.005 383.405 ;
      END
   END dout1[54]
   PIN dout1[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  519.865 383.025 520.245 383.405 ;
      END
   END dout1[55]
   PIN dout1[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  526.105 383.025 526.485 383.405 ;
      END
   END dout1[56]
   PIN dout1[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  532.345 383.025 532.725 383.405 ;
      END
   END dout1[57]
   PIN dout1[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  538.585 383.025 538.965 383.405 ;
      END
   END dout1[58]
   PIN dout1[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  544.825 383.025 545.205 383.405 ;
      END
   END dout1[59]
   PIN dout1[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  551.065 383.025 551.445 383.405 ;
      END
   END dout1[60]
   PIN dout1[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  557.305 383.025 557.685 383.405 ;
      END
   END dout1[61]
   PIN dout1[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  563.545 383.025 563.925 383.405 ;
      END
   END dout1[62]
   PIN dout1[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  569.785 383.025 570.165 383.405 ;
      END
   END dout1[63]
   PIN dout1[64]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  576.025 383.025 576.405 383.405 ;
      END
   END dout1[64]
   PIN dout1[65]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  582.265 383.025 582.645 383.405 ;
      END
   END dout1[65]
   PIN dout1[66]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  588.505 383.025 588.885 383.405 ;
      END
   END dout1[66]
   PIN dout1[67]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  594.745 383.025 595.125 383.405 ;
      END
   END dout1[67]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  0.0 0.0 777.18 1.74 ;
         LAYER met4 ;
         RECT  775.44 0.0 777.18 383.405 ;
         LAYER met3 ;
         RECT  0.0 381.665 777.18 383.405 ;
         LAYER met4 ;
         RECT  0.0 0.0 1.74 383.405 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  771.96 3.48 773.7 379.925 ;
         LAYER met3 ;
         RECT  3.48 3.48 773.7 5.22 ;
         LAYER met4 ;
         RECT  3.48 3.48 5.22 379.925 ;
         LAYER met3 ;
         RECT  3.48 378.185 773.7 379.925 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 776.56 382.785 ;
   LAYER  met2 ;
      RECT  0.62 0.62 776.56 382.785 ;
   LAYER  met3 ;
      RECT  0.98 112.905 776.56 114.485 ;
      RECT  0.62 114.485 0.98 121.405 ;
      RECT  0.62 122.985 0.98 127.275 ;
      RECT  0.62 128.855 0.98 135.675 ;
      RECT  0.62 137.255 0.98 141.185 ;
      RECT  0.62 142.765 0.98 149.685 ;
      RECT  0.62 151.265 0.98 155.325 ;
      RECT  0.62 20.675 0.98 112.905 ;
      RECT  0.98 114.485 776.2 367.555 ;
      RECT  0.98 367.555 776.2 369.135 ;
      RECT  776.2 114.485 776.56 367.555 ;
      RECT  0.62 2.34 0.98 19.095 ;
      RECT  0.62 156.905 0.98 381.065 ;
      RECT  776.2 369.135 776.56 381.065 ;
      RECT  0.98 2.34 2.88 2.88 ;
      RECT  0.98 2.88 2.88 5.82 ;
      RECT  0.98 5.82 2.88 112.905 ;
      RECT  2.88 2.34 774.3 2.88 ;
      RECT  2.88 5.82 774.3 112.905 ;
      RECT  774.3 2.34 776.56 2.88 ;
      RECT  774.3 2.88 776.56 5.82 ;
      RECT  774.3 5.82 776.56 112.905 ;
      RECT  0.98 369.135 2.88 377.585 ;
      RECT  0.98 377.585 2.88 380.525 ;
      RECT  0.98 380.525 2.88 381.065 ;
      RECT  2.88 369.135 774.3 377.585 ;
      RECT  2.88 380.525 774.3 381.065 ;
      RECT  774.3 369.135 776.2 377.585 ;
      RECT  774.3 377.585 776.2 380.525 ;
      RECT  774.3 380.525 776.2 381.065 ;
   LAYER  met4 ;
      RECT  113.34 0.98 114.92 382.785 ;
      RECT  114.92 0.62 119.18 0.98 ;
      RECT  120.76 0.62 125.02 0.98 ;
      RECT  126.6 0.62 130.86 0.98 ;
      RECT  132.44 0.62 136.7 0.98 ;
      RECT  138.28 0.62 142.54 0.98 ;
      RECT  144.12 0.62 148.38 0.98 ;
      RECT  149.96 0.62 154.22 0.98 ;
      RECT  155.8 0.62 160.06 0.98 ;
      RECT  161.64 0.62 165.9 0.98 ;
      RECT  167.48 0.62 171.74 0.98 ;
      RECT  173.32 0.62 177.58 0.98 ;
      RECT  179.16 0.62 183.42 0.98 ;
      RECT  185.0 0.62 189.26 0.98 ;
      RECT  190.84 0.62 195.1 0.98 ;
      RECT  196.68 0.62 200.94 0.98 ;
      RECT  202.52 0.62 206.78 0.98 ;
      RECT  208.36 0.62 212.62 0.98 ;
      RECT  214.2 0.62 218.46 0.98 ;
      RECT  220.04 0.62 224.3 0.98 ;
      RECT  225.88 0.62 230.14 0.98 ;
      RECT  231.72 0.62 235.98 0.98 ;
      RECT  237.56 0.62 241.82 0.98 ;
      RECT  243.4 0.62 247.66 0.98 ;
      RECT  249.24 0.62 253.5 0.98 ;
      RECT  255.08 0.62 259.34 0.98 ;
      RECT  260.92 0.62 265.18 0.98 ;
      RECT  266.76 0.62 271.02 0.98 ;
      RECT  272.6 0.62 276.86 0.98 ;
      RECT  278.44 0.62 282.7 0.98 ;
      RECT  284.28 0.62 288.54 0.98 ;
      RECT  290.12 0.62 294.38 0.98 ;
      RECT  295.96 0.62 300.22 0.98 ;
      RECT  301.8 0.62 306.06 0.98 ;
      RECT  307.64 0.62 311.9 0.98 ;
      RECT  313.48 0.62 317.74 0.98 ;
      RECT  319.32 0.62 323.58 0.98 ;
      RECT  325.16 0.62 329.42 0.98 ;
      RECT  331.0 0.62 335.26 0.98 ;
      RECT  336.84 0.62 341.1 0.98 ;
      RECT  342.68 0.62 346.94 0.98 ;
      RECT  348.52 0.62 352.78 0.98 ;
      RECT  354.36 0.62 358.62 0.98 ;
      RECT  360.2 0.62 364.46 0.98 ;
      RECT  366.04 0.62 370.3 0.98 ;
      RECT  371.88 0.62 376.14 0.98 ;
      RECT  377.72 0.62 381.98 0.98 ;
      RECT  383.56 0.62 387.82 0.98 ;
      RECT  389.4 0.62 393.66 0.98 ;
      RECT  395.24 0.62 399.5 0.98 ;
      RECT  401.08 0.62 405.34 0.98 ;
      RECT  406.92 0.62 411.18 0.98 ;
      RECT  412.76 0.62 417.02 0.98 ;
      RECT  418.6 0.62 422.86 0.98 ;
      RECT  424.44 0.62 428.7 0.98 ;
      RECT  430.28 0.62 434.54 0.98 ;
      RECT  436.12 0.62 440.38 0.98 ;
      RECT  441.96 0.62 446.22 0.98 ;
      RECT  447.8 0.62 452.06 0.98 ;
      RECT  453.64 0.62 457.9 0.98 ;
      RECT  459.48 0.62 463.74 0.98 ;
      RECT  465.32 0.62 469.58 0.98 ;
      RECT  471.16 0.62 475.42 0.98 ;
      RECT  477.0 0.62 481.26 0.98 ;
      RECT  482.84 0.62 487.1 0.98 ;
      RECT  488.68 0.62 492.94 0.98 ;
      RECT  494.52 0.62 498.78 0.98 ;
      RECT  500.36 0.62 504.62 0.98 ;
      RECT  109.08 0.62 113.34 0.98 ;
      RECT  114.92 0.98 662.26 382.425 ;
      RECT  662.26 0.98 663.84 382.425 ;
      RECT  506.2 0.62 676.965 0.98 ;
      RECT  31.24 0.62 107.5 0.98 ;
      RECT  663.84 382.425 745.94 382.785 ;
      RECT  114.92 382.425 176.065 382.785 ;
      RECT  177.645 382.425 182.305 382.785 ;
      RECT  183.885 382.425 188.545 382.785 ;
      RECT  190.125 382.425 194.785 382.785 ;
      RECT  196.365 382.425 201.025 382.785 ;
      RECT  202.605 382.425 207.265 382.785 ;
      RECT  208.845 382.425 213.505 382.785 ;
      RECT  215.085 382.425 219.745 382.785 ;
      RECT  221.325 382.425 225.985 382.785 ;
      RECT  227.565 382.425 232.225 382.785 ;
      RECT  233.805 382.425 238.465 382.785 ;
      RECT  240.045 382.425 244.705 382.785 ;
      RECT  246.285 382.425 250.945 382.785 ;
      RECT  252.525 382.425 257.185 382.785 ;
      RECT  258.765 382.425 263.425 382.785 ;
      RECT  265.005 382.425 269.665 382.785 ;
      RECT  271.245 382.425 275.905 382.785 ;
      RECT  277.485 382.425 282.145 382.785 ;
      RECT  283.725 382.425 288.385 382.785 ;
      RECT  289.965 382.425 294.625 382.785 ;
      RECT  296.205 382.425 300.865 382.785 ;
      RECT  302.445 382.425 307.105 382.785 ;
      RECT  308.685 382.425 313.345 382.785 ;
      RECT  314.925 382.425 319.585 382.785 ;
      RECT  321.165 382.425 325.825 382.785 ;
      RECT  327.405 382.425 332.065 382.785 ;
      RECT  333.645 382.425 338.305 382.785 ;
      RECT  339.885 382.425 344.545 382.785 ;
      RECT  346.125 382.425 350.785 382.785 ;
      RECT  352.365 382.425 357.025 382.785 ;
      RECT  358.605 382.425 363.265 382.785 ;
      RECT  364.845 382.425 369.505 382.785 ;
      RECT  371.085 382.425 375.745 382.785 ;
      RECT  377.325 382.425 381.985 382.785 ;
      RECT  383.565 382.425 388.225 382.785 ;
      RECT  389.805 382.425 394.465 382.785 ;
      RECT  396.045 382.425 400.705 382.785 ;
      RECT  402.285 382.425 406.945 382.785 ;
      RECT  408.525 382.425 413.185 382.785 ;
      RECT  414.765 382.425 419.425 382.785 ;
      RECT  421.005 382.425 425.665 382.785 ;
      RECT  427.245 382.425 431.905 382.785 ;
      RECT  433.485 382.425 438.145 382.785 ;
      RECT  439.725 382.425 444.385 382.785 ;
      RECT  445.965 382.425 450.625 382.785 ;
      RECT  452.205 382.425 456.865 382.785 ;
      RECT  458.445 382.425 463.105 382.785 ;
      RECT  464.685 382.425 469.345 382.785 ;
      RECT  470.925 382.425 475.585 382.785 ;
      RECT  477.165 382.425 481.825 382.785 ;
      RECT  483.405 382.425 488.065 382.785 ;
      RECT  489.645 382.425 494.305 382.785 ;
      RECT  495.885 382.425 500.545 382.785 ;
      RECT  502.125 382.425 506.785 382.785 ;
      RECT  508.365 382.425 513.025 382.785 ;
      RECT  514.605 382.425 519.265 382.785 ;
      RECT  520.845 382.425 525.505 382.785 ;
      RECT  527.085 382.425 531.745 382.785 ;
      RECT  533.325 382.425 537.985 382.785 ;
      RECT  539.565 382.425 544.225 382.785 ;
      RECT  545.805 382.425 550.465 382.785 ;
      RECT  552.045 382.425 556.705 382.785 ;
      RECT  558.285 382.425 562.945 382.785 ;
      RECT  564.525 382.425 569.185 382.785 ;
      RECT  570.765 382.425 575.425 382.785 ;
      RECT  577.005 382.425 581.665 382.785 ;
      RECT  583.245 382.425 587.905 382.785 ;
      RECT  589.485 382.425 594.145 382.785 ;
      RECT  595.725 382.425 662.26 382.785 ;
      RECT  683.59 0.62 774.84 0.98 ;
      RECT  747.52 382.425 774.84 382.785 ;
      RECT  2.34 0.62 29.66 0.98 ;
      RECT  663.84 0.98 771.36 2.88 ;
      RECT  663.84 2.88 771.36 380.525 ;
      RECT  663.84 380.525 771.36 382.425 ;
      RECT  771.36 0.98 774.3 2.88 ;
      RECT  771.36 380.525 774.3 382.425 ;
      RECT  774.3 0.98 774.84 2.88 ;
      RECT  774.3 2.88 774.84 380.525 ;
      RECT  774.3 380.525 774.84 382.425 ;
      RECT  2.34 0.98 2.88 2.88 ;
      RECT  2.34 2.88 2.88 380.525 ;
      RECT  2.34 380.525 2.88 382.785 ;
      RECT  2.88 0.98 5.82 2.88 ;
      RECT  2.88 380.525 5.82 382.785 ;
      RECT  5.82 0.98 113.34 2.88 ;
      RECT  5.82 2.88 113.34 380.525 ;
      RECT  5.82 380.525 113.34 382.785 ;
   END
END    sky130_sram_1r1w0rw_68x256
END    LIBRARY
